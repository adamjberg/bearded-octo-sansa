// nios_system.v

// Generated using ACDS version 12.0sp2 263 at 2013.02.16.18:56:48

`timescale 1 ps / 1 ps
module nios_system (
		output wire        vga_extern_CLK,                          //                         vga_extern.CLK
		output wire        vga_extern_HS,                           //                                   .HS
		output wire        vga_extern_VS,                           //                                   .VS
		output wire        vga_extern_BLANK,                        //                                   .BLANK
		output wire        vga_extern_SYNC,                         //                                   .SYNC
		output wire [9:0]  vga_extern_R,                            //                                   .R
		output wire [9:0]  vga_extern_G,                            //                                   .G
		output wire [9:0]  vga_extern_B,                            //                                   .B
		input  wire        clk_in_secondary_clk,                    //                   clk_in_secondary.clk
		input  wire        audio_ADCDAT,                            //                              audio.ADCDAT
		input  wire        audio_ADCLRCK,                           //                                   .ADCLRCK
		input  wire        audio_BCLK,                              //                                   .BCLK
		output wire        audio_DACDAT,                            //                                   .DACDAT
		input  wire        audio_DACLRCK,                           //                                   .DACLRCK
		inout  wire        sd_card_b_SD_cmd,                        //                            sd_card.b_SD_cmd
		inout  wire        sd_card_b_SD_dat,                        //                                   .b_SD_dat
		inout  wire        sd_card_b_SD_dat3,                       //                                   .b_SD_dat3
		output wire        sd_card_o_SD_clock,                      //                                   .o_SD_clock
		input  wire [3:0]  keys_export,                             //                               keys.export
		input  wire        clk_clk,                                 //                                clk.clk
		output wire [7:0]  hex2_ex_export,                          //                            hex2_ex.export
		inout  wire        ps2_0_external_interface_CLK,            //           ps2_0_external_interface.CLK
		inout  wire        ps2_0_external_interface_DAT,            //                                   .DAT
		output wire        audio_clk_clk,                           //                          audio_clk.clk
		inout  wire [15:0] sram_interface_DQ,                       //                     sram_interface.DQ
		output wire [17:0] sram_interface_ADDR,                     //                                   .ADDR
		output wire        sram_interface_LB_N,                     //                                   .LB_N
		output wire        sram_interface_UB_N,                     //                                   .UB_N
		output wire        sram_interface_CE_N,                     //                                   .CE_N
		output wire        sram_interface_OE_N,                     //                                   .OE_N
		output wire        sram_interface_WE_N,                     //                                   .WE_N
		input  wire [7:0]  switches_export,                         //                           switches.export
		output wire [17:0] ledrs_export,                            //                              ledrs.export
		output wire [7:0]  hex0_ex_export,                          //                            hex0_ex.export
		output wire [7:0]  leds_export,                             //                               leds.export
		inout  wire [7:0]  character_lcd_0_external_interface_DATA, // character_lcd_0_external_interface.DATA
		output wire        character_lcd_0_external_interface_ON,   //                                   .ON
		output wire        character_lcd_0_external_interface_BLON, //                                   .BLON
		output wire        character_lcd_0_external_interface_EN,   //                                   .EN
		output wire        character_lcd_0_external_interface_RS,   //                                   .RS
		output wire        character_lcd_0_external_interface_RW,   //                                   .RW
		output wire [7:0]  hex3_ex_export,                          //                            hex3_ex.export
		output wire [11:0] sdram_wire_addr,                         //                         sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                           //                                   .ba
		output wire        sdram_wire_cas_n,                        //                                   .cas_n
		output wire        sdram_wire_cke,                          //                                   .cke
		output wire        sdram_wire_cs_n,                         //                                   .cs_n
		inout  wire [15:0] sdram_wire_dq,                           //                                   .dq
		output wire [1:0]  sdram_wire_dqm,                          //                                   .dqm
		output wire        sdram_wire_ras_n,                        //                                   .ras_n
		output wire        sdram_wire_we_n,                         //                                   .we_n
		input  wire        reset_reset_n,                           //                              reset.reset_n
		output wire [7:0]  hex1_ex_export,                          //                            hex1_ex.export
		output wire [7:0]  hex4_ex_export,                          //                            hex4_ex.export
		inout  wire        audio_and_video_config_SDAT,             //             audio_and_video_config.SDAT
		output wire        audio_and_video_config_SCLK,             //                                   .SCLK
		output wire        sdram_clk_clk                            //                          sdram_clk.clk
	);

	wire          clocks_sys_clk_clk;                                                                                                   // clocks:sys_clk -> [Keys:clk, Keys_s1_translator:clk, Keys_s1_translator_avalon_universal_slave_0_agent:clk, Keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, LEDR:clk, LEDR_s1_translator:clk, LEDR_s1_translator_avalon_universal_slave_0_agent:clk, LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, SD_Card:i_clock, SD_Card_avalon_sdcard_slave_translator:clk, SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:clk, SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Switches:clk, Switches_s1_translator:clk, Switches_s1_translator_avalon_universal_slave_0_agent:clk, Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, addr_router_001:clk, addr_router_002:clk, alpha_blender:clk, audio:clk, audio_and_video_config_0:clk, audio_and_video_config_0_avalon_av_config_slave_translator:clk, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:clk, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, audio_avalon_audio_slave_translator:clk, audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:clk, audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, burst_adapter:clk, burst_adapter_001:clk, burst_adapter_002:clk, burst_adapter_003:clk, char_drawer:clk, char_drawer_avalon_char_buffer_slave_translator:clk, char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:clk, char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, char_drawer_avalon_char_control_slave_translator:clk, char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:clk, char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, character_lcd_0:clk, character_lcd_0_avalon_lcd_slave_translator:clk, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:clk, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_005:clk, hex0:clk, hex0_s1_translator:clk, hex0_s1_translator_avalon_universal_slave_0_agent:clk, hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, hex1:clk, hex1_s1_translator:clk, hex1_s1_translator_avalon_universal_slave_0_agent:clk, hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, hex2:clk, hex2_s1_translator:clk, hex2_s1_translator_avalon_universal_slave_0_agent:clk, hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, hex3:clk, hex3_s1_translator:clk, hex3_s1_translator_avalon_universal_slave_0_agent:clk, hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, hex4:clk, hex4_s1_translator:clk, hex4_s1_translator_avalon_universal_slave_0_agent:clk, hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, id_router_016:clk, id_router_017:clk, id_router_018:clk, id_router_019:clk, id_router_020:clk, id_router_021:clk, id_router_022:clk, irq_mapper:clk, jtag_uart:clk, jtag_uart_avalon_jtag_slave_translator:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, leds:clk, leds_s1_translator:clk, leds_s1_translator_avalon_universal_slave_0_agent:clk, leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter:clk, limiter_001:clk, nios2_processor:clk, nios2_processor_data_master_translator:clk, nios2_processor_data_master_translator_avalon_universal_master_0_agent:clk, nios2_processor_instruction_master_translator:clk, nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_processor_jtag_debug_module_translator:clk, nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pixel_buffer:clk, pixel_buffer_avalon_sram_slave_translator:clk, pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pixel_buffer_dma_0:clk, pixel_buffer_dma_0_avalon_control_slave_translator:clk, pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:clk, pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pixel_buffer_dma_0_avalon_pixel_dma_master_translator:clk, pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:clk, ps2_0:clk, ps2_0_avalon_ps2_slave_translator:clk, ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:clk, ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rgb_resampler:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_demux_016:clk, rsp_xbar_demux_017:clk, rsp_xbar_demux_018:clk, rsp_xbar_demux_019:clk, rsp_xbar_demux_020:clk, rsp_xbar_demux_021:clk, rsp_xbar_demux_022:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, rst_controller_003:clk, scaler:clk, sdram:clk, sdram_s1_translator:clk, sdram_s1_translator_avalon_universal_slave_0_agent:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer:clk, timer_s1_translator:clk, timer_s1_translator_avalon_universal_slave_0_agent:clk, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timestamp:clk, timestamp_s1_translator:clk, timestamp_s1_translator_avalon_universal_slave_0_agent:clk, timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, up_clocks_0:CLOCK_50, video_fifo:clk_stream_in, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk, width_adapter_006:clk, width_adapter_007:clk, width_adapter_008:clk, width_adapter_009:clk]
	wire          pixel_buffer_dma_0_avalon_pixel_source_endofpacket;                                                                   // pixel_buffer_dma_0:stream_endofpacket -> rgb_resampler:stream_in_endofpacket
	wire          pixel_buffer_dma_0_avalon_pixel_source_valid;                                                                         // pixel_buffer_dma_0:stream_valid -> rgb_resampler:stream_in_valid
	wire          pixel_buffer_dma_0_avalon_pixel_source_startofpacket;                                                                 // pixel_buffer_dma_0:stream_startofpacket -> rgb_resampler:stream_in_startofpacket
	wire   [15:0] pixel_buffer_dma_0_avalon_pixel_source_data;                                                                          // pixel_buffer_dma_0:stream_data -> rgb_resampler:stream_in_data
	wire          pixel_buffer_dma_0_avalon_pixel_source_ready;                                                                         // rgb_resampler:stream_in_ready -> pixel_buffer_dma_0:stream_ready
	wire          rgb_resampler_avalon_rgb_source_endofpacket;                                                                          // rgb_resampler:stream_out_endofpacket -> scaler:stream_in_endofpacket
	wire          rgb_resampler_avalon_rgb_source_valid;                                                                                // rgb_resampler:stream_out_valid -> scaler:stream_in_valid
	wire          rgb_resampler_avalon_rgb_source_startofpacket;                                                                        // rgb_resampler:stream_out_startofpacket -> scaler:stream_in_startofpacket
	wire   [29:0] rgb_resampler_avalon_rgb_source_data;                                                                                 // rgb_resampler:stream_out_data -> scaler:stream_in_data
	wire          rgb_resampler_avalon_rgb_source_ready;                                                                                // scaler:stream_in_ready -> rgb_resampler:stream_out_ready
	wire          video_fifo_avalon_dc_buffer_source_endofpacket;                                                                       // video_fifo:stream_out_endofpacket -> vga_controller:endofpacket
	wire          video_fifo_avalon_dc_buffer_source_valid;                                                                             // video_fifo:stream_out_valid -> vga_controller:valid
	wire          video_fifo_avalon_dc_buffer_source_startofpacket;                                                                     // video_fifo:stream_out_startofpacket -> vga_controller:startofpacket
	wire   [29:0] video_fifo_avalon_dc_buffer_source_data;                                                                              // video_fifo:stream_out_data -> vga_controller:data
	wire          video_fifo_avalon_dc_buffer_source_ready;                                                                             // vga_controller:ready -> video_fifo:stream_out_ready
	wire          char_drawer_avalon_char_source_endofpacket;                                                                           // char_drawer:stream_endofpacket -> alpha_blender:foreground_endofpacket
	wire          char_drawer_avalon_char_source_valid;                                                                                 // char_drawer:stream_valid -> alpha_blender:foreground_valid
	wire          char_drawer_avalon_char_source_startofpacket;                                                                         // char_drawer:stream_startofpacket -> alpha_blender:foreground_startofpacket
	wire   [39:0] char_drawer_avalon_char_source_data;                                                                                  // char_drawer:stream_data -> alpha_blender:foreground_data
	wire          char_drawer_avalon_char_source_ready;                                                                                 // alpha_blender:foreground_ready -> char_drawer:stream_ready
	wire          scaler_avalon_scaler_source_endofpacket;                                                                              // scaler:stream_out_endofpacket -> alpha_blender:background_endofpacket
	wire          scaler_avalon_scaler_source_valid;                                                                                    // scaler:stream_out_valid -> alpha_blender:background_valid
	wire          scaler_avalon_scaler_source_startofpacket;                                                                            // scaler:stream_out_startofpacket -> alpha_blender:background_startofpacket
	wire   [29:0] scaler_avalon_scaler_source_data;                                                                                     // scaler:stream_out_data -> alpha_blender:background_data
	wire          scaler_avalon_scaler_source_ready;                                                                                    // alpha_blender:background_ready -> scaler:stream_out_ready
	wire          alpha_blender_avalon_blended_source_endofpacket;                                                                      // alpha_blender:output_endofpacket -> video_fifo:stream_in_endofpacket
	wire          alpha_blender_avalon_blended_source_valid;                                                                            // alpha_blender:output_valid -> video_fifo:stream_in_valid
	wire          alpha_blender_avalon_blended_source_startofpacket;                                                                    // alpha_blender:output_startofpacket -> video_fifo:stream_in_startofpacket
	wire   [29:0] alpha_blender_avalon_blended_source_data;                                                                             // alpha_blender:output_data -> video_fifo:stream_in_data
	wire          alpha_blender_avalon_blended_source_ready;                                                                            // video_fifo:stream_in_ready -> alpha_blender:output_ready
	wire          clocks_vga_clk_clk;                                                                                                   // clocks:VGA_CLK -> [rst_controller_002:clk, vga_controller:clk, video_fifo:clk_stream_out]
	wire          nios2_processor_instruction_master_waitrequest;                                                                       // nios2_processor_instruction_master_translator:av_waitrequest -> nios2_processor:i_waitrequest
	wire   [24:0] nios2_processor_instruction_master_address;                                                                           // nios2_processor:i_address -> nios2_processor_instruction_master_translator:av_address
	wire          nios2_processor_instruction_master_read;                                                                              // nios2_processor:i_read -> nios2_processor_instruction_master_translator:av_read
	wire   [31:0] nios2_processor_instruction_master_readdata;                                                                          // nios2_processor_instruction_master_translator:av_readdata -> nios2_processor:i_readdata
	wire          nios2_processor_instruction_master_readdatavalid;                                                                     // nios2_processor_instruction_master_translator:av_readdatavalid -> nios2_processor:i_readdatavalid
	wire          nios2_processor_data_master_waitrequest;                                                                              // nios2_processor_data_master_translator:av_waitrequest -> nios2_processor:d_waitrequest
	wire   [31:0] nios2_processor_data_master_writedata;                                                                                // nios2_processor:d_writedata -> nios2_processor_data_master_translator:av_writedata
	wire   [24:0] nios2_processor_data_master_address;                                                                                  // nios2_processor:d_address -> nios2_processor_data_master_translator:av_address
	wire          nios2_processor_data_master_write;                                                                                    // nios2_processor:d_write -> nios2_processor_data_master_translator:av_write
	wire          nios2_processor_data_master_read;                                                                                     // nios2_processor:d_read -> nios2_processor_data_master_translator:av_read
	wire   [31:0] nios2_processor_data_master_readdata;                                                                                 // nios2_processor_data_master_translator:av_readdata -> nios2_processor:d_readdata
	wire          nios2_processor_data_master_debugaccess;                                                                              // nios2_processor:jtag_debug_module_debugaccess_to_roms -> nios2_processor_data_master_translator:av_debugaccess
	wire          nios2_processor_data_master_readdatavalid;                                                                            // nios2_processor_data_master_translator:av_readdatavalid -> nios2_processor:d_readdatavalid
	wire    [3:0] nios2_processor_data_master_byteenable;                                                                               // nios2_processor:d_byteenable -> nios2_processor_data_master_translator:av_byteenable
	wire          pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest;                                                               // pixel_buffer_dma_0_avalon_pixel_dma_master_translator:av_waitrequest -> pixel_buffer_dma_0:master_waitrequest
	wire   [31:0] pixel_buffer_dma_0_avalon_pixel_dma_master_address;                                                                   // pixel_buffer_dma_0:master_address -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator:av_address
	wire          pixel_buffer_dma_0_avalon_pixel_dma_master_lock;                                                                      // pixel_buffer_dma_0:master_arbiterlock -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator:av_lock
	wire          pixel_buffer_dma_0_avalon_pixel_dma_master_read;                                                                      // pixel_buffer_dma_0:master_read -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator:av_read
	wire   [15:0] pixel_buffer_dma_0_avalon_pixel_dma_master_readdata;                                                                  // pixel_buffer_dma_0_avalon_pixel_dma_master_translator:av_readdata -> pixel_buffer_dma_0:master_readdata
	wire          pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid;                                                             // pixel_buffer_dma_0_avalon_pixel_dma_master_translator:av_readdatavalid -> pixel_buffer_dma_0:master_readdatavalid
	wire   [31:0] nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                           // nios2_processor_jtag_debug_module_translator:av_writedata -> nios2_processor:jtag_debug_module_writedata
	wire    [8:0] nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_address;                                             // nios2_processor_jtag_debug_module_translator:av_address -> nios2_processor:jtag_debug_module_address
	wire          nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                          // nios2_processor_jtag_debug_module_translator:av_chipselect -> nios2_processor:jtag_debug_module_select
	wire          nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_write;                                               // nios2_processor_jtag_debug_module_translator:av_write -> nios2_processor:jtag_debug_module_write
	wire   [31:0] nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                            // nios2_processor:jtag_debug_module_readdata -> nios2_processor_jtag_debug_module_translator:av_readdata
	wire          nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                       // nios2_processor_jtag_debug_module_translator:av_begintransfer -> nios2_processor:jtag_debug_module_begintransfer
	wire          nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                         // nios2_processor_jtag_debug_module_translator:av_debugaccess -> nios2_processor:jtag_debug_module_debugaccess
	wire    [3:0] nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                          // nios2_processor_jtag_debug_module_translator:av_byteenable -> nios2_processor:jtag_debug_module_byteenable
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                                                  // sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                                    // sdram_s1_translator:av_writedata -> sdram:az_data
	wire   [21:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                                      // sdram_s1_translator:av_address -> sdram:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                                                   // sdram_s1_translator:av_chipselect -> sdram:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                                        // sdram_s1_translator:av_write -> sdram:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                                         // sdram_s1_translator:av_read -> sdram:az_rd_n
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                                     // sdram:za_data -> sdram_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                                                // sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	wire    [1:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                                                   // sdram_s1_translator:av_byteenable -> sdram:az_be_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                               // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                                 // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                                   // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                                // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                                     // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                                      // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                                  // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_writedata;                                                                    // timer_s1_translator:av_writedata -> timer:writedata
	wire    [2:0] timer_s1_translator_avalon_anti_slave_0_address;                                                                      // timer_s1_translator:av_address -> timer:address
	wire          timer_s1_translator_avalon_anti_slave_0_chipselect;                                                                   // timer_s1_translator:av_chipselect -> timer:chipselect
	wire          timer_s1_translator_avalon_anti_slave_0_write;                                                                        // timer_s1_translator:av_write -> timer:write_n
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_readdata;                                                                     // timer:readdata -> timer_s1_translator:av_readdata
	wire   [15:0] timestamp_s1_translator_avalon_anti_slave_0_writedata;                                                                // timestamp_s1_translator:av_writedata -> timestamp:writedata
	wire    [2:0] timestamp_s1_translator_avalon_anti_slave_0_address;                                                                  // timestamp_s1_translator:av_address -> timestamp:address
	wire          timestamp_s1_translator_avalon_anti_slave_0_chipselect;                                                               // timestamp_s1_translator:av_chipselect -> timestamp:chipselect
	wire          timestamp_s1_translator_avalon_anti_slave_0_write;                                                                    // timestamp_s1_translator:av_write -> timestamp:write_n
	wire   [15:0] timestamp_s1_translator_avalon_anti_slave_0_readdata;                                                                 // timestamp:readdata -> timestamp_s1_translator:av_readdata
	wire   [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata;                                              // pixel_buffer_avalon_sram_slave_translator:av_writedata -> pixel_buffer:writedata
	wire   [17:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address;                                                // pixel_buffer_avalon_sram_slave_translator:av_address -> pixel_buffer:address
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write;                                                  // pixel_buffer_avalon_sram_slave_translator:av_write -> pixel_buffer:write
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read;                                                   // pixel_buffer_avalon_sram_slave_translator:av_read -> pixel_buffer:read
	wire   [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata;                                               // pixel_buffer:readdata -> pixel_buffer_avalon_sram_slave_translator:av_readdata
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid;                                          // pixel_buffer:readdatavalid -> pixel_buffer_avalon_sram_slave_translator:av_readdatavalid
	wire    [1:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable;                                             // pixel_buffer_avalon_sram_slave_translator:av_byteenable -> pixel_buffer:byteenable
	wire   [31:0] pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_writedata;                                     // pixel_buffer_dma_0_avalon_control_slave_translator:av_writedata -> pixel_buffer_dma_0:slave_writedata
	wire    [1:0] pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_address;                                       // pixel_buffer_dma_0_avalon_control_slave_translator:av_address -> pixel_buffer_dma_0:slave_address
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_write;                                         // pixel_buffer_dma_0_avalon_control_slave_translator:av_write -> pixel_buffer_dma_0:slave_write
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_read;                                          // pixel_buffer_dma_0_avalon_control_slave_translator:av_read -> pixel_buffer_dma_0:slave_read
	wire   [31:0] pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_readdata;                                      // pixel_buffer_dma_0:slave_readdata -> pixel_buffer_dma_0_avalon_control_slave_translator:av_readdata
	wire    [3:0] pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_byteenable;                                    // pixel_buffer_dma_0_avalon_control_slave_translator:av_byteenable -> pixel_buffer_dma_0:slave_byteenable
	wire   [31:0] char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata;                                       // char_drawer_avalon_char_control_slave_translator:av_writedata -> char_drawer:ctrl_writedata
	wire          char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_address;                                         // char_drawer_avalon_char_control_slave_translator:av_address -> char_drawer:ctrl_address
	wire          char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect;                                      // char_drawer_avalon_char_control_slave_translator:av_chipselect -> char_drawer:ctrl_chipselect
	wire          char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_write;                                           // char_drawer_avalon_char_control_slave_translator:av_write -> char_drawer:ctrl_write
	wire          char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_read;                                            // char_drawer_avalon_char_control_slave_translator:av_read -> char_drawer:ctrl_read
	wire   [31:0] char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata;                                        // char_drawer:ctrl_readdata -> char_drawer_avalon_char_control_slave_translator:av_readdata
	wire    [3:0] char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable;                                      // char_drawer_avalon_char_control_slave_translator:av_byteenable -> char_drawer:ctrl_byteenable
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest;                                      // char_drawer:buf_waitrequest -> char_drawer_avalon_char_buffer_slave_translator:av_waitrequest
	wire    [7:0] char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata;                                        // char_drawer_avalon_char_buffer_slave_translator:av_writedata -> char_drawer:buf_writedata
	wire   [12:0] char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address;                                          // char_drawer_avalon_char_buffer_slave_translator:av_address -> char_drawer:buf_address
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect;                                       // char_drawer_avalon_char_buffer_slave_translator:av_chipselect -> char_drawer:buf_chipselect
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write;                                            // char_drawer_avalon_char_buffer_slave_translator:av_write -> char_drawer:buf_write
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read;                                             // char_drawer_avalon_char_buffer_slave_translator:av_read -> char_drawer:buf_read
	wire    [7:0] char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata;                                         // char_drawer:buf_readdata -> char_drawer_avalon_char_buffer_slave_translator:av_readdata
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable;                                       // char_drawer_avalon_char_buffer_slave_translator:av_byteenable -> char_drawer:buf_byteenable
	wire   [31:0] leds_s1_translator_avalon_anti_slave_0_writedata;                                                                     // leds_s1_translator:av_writedata -> leds:writedata
	wire    [1:0] leds_s1_translator_avalon_anti_slave_0_address;                                                                       // leds_s1_translator:av_address -> leds:address
	wire          leds_s1_translator_avalon_anti_slave_0_chipselect;                                                                    // leds_s1_translator:av_chipselect -> leds:chipselect
	wire          leds_s1_translator_avalon_anti_slave_0_write;                                                                         // leds_s1_translator:av_write -> leds:write_n
	wire   [31:0] leds_s1_translator_avalon_anti_slave_0_readdata;                                                                      // leds:readdata -> leds_s1_translator:av_readdata
	wire          sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest;                                               // SD_Card:o_avalon_waitrequest -> SD_Card_avalon_sdcard_slave_translator:av_waitrequest
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata;                                                 // SD_Card_avalon_sdcard_slave_translator:av_writedata -> SD_Card:i_avalon_writedata
	wire    [7:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_address;                                                   // SD_Card_avalon_sdcard_slave_translator:av_address -> SD_Card:i_avalon_address
	wire          sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect;                                                // SD_Card_avalon_sdcard_slave_translator:av_chipselect -> SD_Card:i_avalon_chip_select
	wire          sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_write;                                                     // SD_Card_avalon_sdcard_slave_translator:av_write -> SD_Card:i_avalon_write
	wire          sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_read;                                                      // SD_Card_avalon_sdcard_slave_translator:av_read -> SD_Card:i_avalon_read
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata;                                                  // SD_Card:o_avalon_readdata -> SD_Card_avalon_sdcard_slave_translator:av_readdata
	wire    [3:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable;                                                // SD_Card_avalon_sdcard_slave_translator:av_byteenable -> SD_Card:i_avalon_byteenable
	wire   [31:0] switches_s1_translator_avalon_anti_slave_0_writedata;                                                                 // Switches_s1_translator:av_writedata -> Switches:writedata
	wire    [1:0] switches_s1_translator_avalon_anti_slave_0_address;                                                                   // Switches_s1_translator:av_address -> Switches:address
	wire          switches_s1_translator_avalon_anti_slave_0_chipselect;                                                                // Switches_s1_translator:av_chipselect -> Switches:chipselect
	wire          switches_s1_translator_avalon_anti_slave_0_write;                                                                     // Switches_s1_translator:av_write -> Switches:write_n
	wire   [31:0] switches_s1_translator_avalon_anti_slave_0_readdata;                                                                  // Switches:readdata -> Switches_s1_translator:av_readdata
	wire   [31:0] keys_s1_translator_avalon_anti_slave_0_writedata;                                                                     // Keys_s1_translator:av_writedata -> Keys:writedata
	wire    [1:0] keys_s1_translator_avalon_anti_slave_0_address;                                                                       // Keys_s1_translator:av_address -> Keys:address
	wire          keys_s1_translator_avalon_anti_slave_0_chipselect;                                                                    // Keys_s1_translator:av_chipselect -> Keys:chipselect
	wire          keys_s1_translator_avalon_anti_slave_0_write;                                                                         // Keys_s1_translator:av_write -> Keys:write_n
	wire   [31:0] keys_s1_translator_avalon_anti_slave_0_readdata;                                                                      // Keys:readdata -> Keys_s1_translator:av_readdata
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest;                           // audio_and_video_config_0:waitrequest -> audio_and_video_config_0_avalon_av_config_slave_translator:av_waitrequest
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata;                             // audio_and_video_config_0_avalon_av_config_slave_translator:av_writedata -> audio_and_video_config_0:writedata
	wire    [1:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_address;                               // audio_and_video_config_0_avalon_av_config_slave_translator:av_address -> audio_and_video_config_0:address
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_write;                                 // audio_and_video_config_0_avalon_av_config_slave_translator:av_write -> audio_and_video_config_0:write
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_read;                                  // audio_and_video_config_0_avalon_av_config_slave_translator:av_read -> audio_and_video_config_0:read
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata;                              // audio_and_video_config_0:readdata -> audio_and_video_config_0_avalon_av_config_slave_translator:av_readdata
	wire    [3:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable;                            // audio_and_video_config_0_avalon_av_config_slave_translator:av_byteenable -> audio_and_video_config_0:byteenable
	wire   [31:0] audio_avalon_audio_slave_translator_avalon_anti_slave_0_writedata;                                                    // audio_avalon_audio_slave_translator:av_writedata -> audio:writedata
	wire    [1:0] audio_avalon_audio_slave_translator_avalon_anti_slave_0_address;                                                      // audio_avalon_audio_slave_translator:av_address -> audio:address
	wire          audio_avalon_audio_slave_translator_avalon_anti_slave_0_chipselect;                                                   // audio_avalon_audio_slave_translator:av_chipselect -> audio:chipselect
	wire          audio_avalon_audio_slave_translator_avalon_anti_slave_0_write;                                                        // audio_avalon_audio_slave_translator:av_write -> audio:write
	wire          audio_avalon_audio_slave_translator_avalon_anti_slave_0_read;                                                         // audio_avalon_audio_slave_translator:av_read -> audio:read
	wire   [31:0] audio_avalon_audio_slave_translator_avalon_anti_slave_0_readdata;                                                     // audio:readdata -> audio_avalon_audio_slave_translator:av_readdata
	wire   [31:0] ledr_s1_translator_avalon_anti_slave_0_writedata;                                                                     // LEDR_s1_translator:av_writedata -> LEDR:writedata
	wire    [1:0] ledr_s1_translator_avalon_anti_slave_0_address;                                                                       // LEDR_s1_translator:av_address -> LEDR:address
	wire          ledr_s1_translator_avalon_anti_slave_0_chipselect;                                                                    // LEDR_s1_translator:av_chipselect -> LEDR:chipselect
	wire          ledr_s1_translator_avalon_anti_slave_0_write;                                                                         // LEDR_s1_translator:av_write -> LEDR:write_n
	wire   [31:0] ledr_s1_translator_avalon_anti_slave_0_readdata;                                                                      // LEDR:readdata -> LEDR_s1_translator:av_readdata
	wire          ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_waitrequest;                                                    // ps2_0:waitrequest -> ps2_0_avalon_ps2_slave_translator:av_waitrequest
	wire   [31:0] ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_writedata;                                                      // ps2_0_avalon_ps2_slave_translator:av_writedata -> ps2_0:writedata
	wire          ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_address;                                                        // ps2_0_avalon_ps2_slave_translator:av_address -> ps2_0:address
	wire          ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_chipselect;                                                     // ps2_0_avalon_ps2_slave_translator:av_chipselect -> ps2_0:chipselect
	wire          ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_write;                                                          // ps2_0_avalon_ps2_slave_translator:av_write -> ps2_0:write
	wire          ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_read;                                                           // ps2_0_avalon_ps2_slave_translator:av_read -> ps2_0:read
	wire   [31:0] ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_readdata;                                                       // ps2_0:readdata -> ps2_0_avalon_ps2_slave_translator:av_readdata
	wire    [3:0] ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_byteenable;                                                     // ps2_0_avalon_ps2_slave_translator:av_byteenable -> ps2_0:byteenable
	wire   [31:0] hex0_s1_translator_avalon_anti_slave_0_writedata;                                                                     // hex0_s1_translator:av_writedata -> hex0:writedata
	wire    [1:0] hex0_s1_translator_avalon_anti_slave_0_address;                                                                       // hex0_s1_translator:av_address -> hex0:address
	wire          hex0_s1_translator_avalon_anti_slave_0_chipselect;                                                                    // hex0_s1_translator:av_chipselect -> hex0:chipselect
	wire          hex0_s1_translator_avalon_anti_slave_0_write;                                                                         // hex0_s1_translator:av_write -> hex0:write_n
	wire   [31:0] hex0_s1_translator_avalon_anti_slave_0_readdata;                                                                      // hex0:readdata -> hex0_s1_translator:av_readdata
	wire   [31:0] hex1_s1_translator_avalon_anti_slave_0_writedata;                                                                     // hex1_s1_translator:av_writedata -> hex1:writedata
	wire    [1:0] hex1_s1_translator_avalon_anti_slave_0_address;                                                                       // hex1_s1_translator:av_address -> hex1:address
	wire          hex1_s1_translator_avalon_anti_slave_0_chipselect;                                                                    // hex1_s1_translator:av_chipselect -> hex1:chipselect
	wire          hex1_s1_translator_avalon_anti_slave_0_write;                                                                         // hex1_s1_translator:av_write -> hex1:write_n
	wire   [31:0] hex1_s1_translator_avalon_anti_slave_0_readdata;                                                                      // hex1:readdata -> hex1_s1_translator:av_readdata
	wire   [31:0] hex2_s1_translator_avalon_anti_slave_0_writedata;                                                                     // hex2_s1_translator:av_writedata -> hex2:writedata
	wire    [1:0] hex2_s1_translator_avalon_anti_slave_0_address;                                                                       // hex2_s1_translator:av_address -> hex2:address
	wire          hex2_s1_translator_avalon_anti_slave_0_chipselect;                                                                    // hex2_s1_translator:av_chipselect -> hex2:chipselect
	wire          hex2_s1_translator_avalon_anti_slave_0_write;                                                                         // hex2_s1_translator:av_write -> hex2:write_n
	wire   [31:0] hex2_s1_translator_avalon_anti_slave_0_readdata;                                                                      // hex2:readdata -> hex2_s1_translator:av_readdata
	wire   [31:0] hex3_s1_translator_avalon_anti_slave_0_writedata;                                                                     // hex3_s1_translator:av_writedata -> hex3:writedata
	wire    [1:0] hex3_s1_translator_avalon_anti_slave_0_address;                                                                       // hex3_s1_translator:av_address -> hex3:address
	wire          hex3_s1_translator_avalon_anti_slave_0_chipselect;                                                                    // hex3_s1_translator:av_chipselect -> hex3:chipselect
	wire          hex3_s1_translator_avalon_anti_slave_0_write;                                                                         // hex3_s1_translator:av_write -> hex3:write_n
	wire   [31:0] hex3_s1_translator_avalon_anti_slave_0_readdata;                                                                      // hex3:readdata -> hex3_s1_translator:av_readdata
	wire   [31:0] hex4_s1_translator_avalon_anti_slave_0_writedata;                                                                     // hex4_s1_translator:av_writedata -> hex4:writedata
	wire    [1:0] hex4_s1_translator_avalon_anti_slave_0_address;                                                                       // hex4_s1_translator:av_address -> hex4:address
	wire          hex4_s1_translator_avalon_anti_slave_0_chipselect;                                                                    // hex4_s1_translator:av_chipselect -> hex4:chipselect
	wire          hex4_s1_translator_avalon_anti_slave_0_write;                                                                         // hex4_s1_translator:av_write -> hex4:write_n
	wire   [31:0] hex4_s1_translator_avalon_anti_slave_0_readdata;                                                                      // hex4:readdata -> hex4_s1_translator:av_readdata
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest;                                          // character_lcd_0:waitrequest -> character_lcd_0_avalon_lcd_slave_translator:av_waitrequest
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata;                                            // character_lcd_0_avalon_lcd_slave_translator:av_writedata -> character_lcd_0:writedata
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address;                                              // character_lcd_0_avalon_lcd_slave_translator:av_address -> character_lcd_0:address
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect;                                           // character_lcd_0_avalon_lcd_slave_translator:av_chipselect -> character_lcd_0:chipselect
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write;                                                // character_lcd_0_avalon_lcd_slave_translator:av_write -> character_lcd_0:write
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read;                                                 // character_lcd_0_avalon_lcd_slave_translator:av_read -> character_lcd_0:read
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata;                                             // character_lcd_0:readdata -> character_lcd_0_avalon_lcd_slave_translator:av_readdata
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_waitrequest;                                  // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_processor_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_burstcount;                                   // nios2_processor_instruction_master_translator:uav_burstcount -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_writedata;                                    // nios2_processor_instruction_master_translator:uav_writedata -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_address;                                      // nios2_processor_instruction_master_translator:uav_address -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_lock;                                         // nios2_processor_instruction_master_translator:uav_lock -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_write;                                        // nios2_processor_instruction_master_translator:uav_write -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_read;                                         // nios2_processor_instruction_master_translator:uav_read -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_readdata;                                     // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_processor_instruction_master_translator:uav_readdata
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_debugaccess;                                  // nios2_processor_instruction_master_translator:uav_debugaccess -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_byteenable;                                   // nios2_processor_instruction_master_translator:uav_byteenable -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_readdatavalid;                                // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_processor_instruction_master_translator:uav_readdatavalid
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_waitrequest;                                         // nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_processor_data_master_translator:uav_waitrequest
	wire    [2:0] nios2_processor_data_master_translator_avalon_universal_master_0_burstcount;                                          // nios2_processor_data_master_translator:uav_burstcount -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_processor_data_master_translator_avalon_universal_master_0_writedata;                                           // nios2_processor_data_master_translator:uav_writedata -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_processor_data_master_translator_avalon_universal_master_0_address;                                             // nios2_processor_data_master_translator:uav_address -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_lock;                                                // nios2_processor_data_master_translator:uav_lock -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_write;                                               // nios2_processor_data_master_translator:uav_write -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_read;                                                // nios2_processor_data_master_translator:uav_read -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_processor_data_master_translator_avalon_universal_master_0_readdata;                                            // nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_processor_data_master_translator:uav_readdata
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_debugaccess;                                         // nios2_processor_data_master_translator:uav_debugaccess -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_processor_data_master_translator_avalon_universal_master_0_byteenable;                                          // nios2_processor_data_master_translator:uav_byteenable -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_readdatavalid;                                       // nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_processor_data_master_translator:uav_readdatavalid
	wire          pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest;                          // pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator:uav_waitrequest
	wire    [1:0] pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount;                           // pixel_buffer_dma_0_avalon_pixel_dma_master_translator:uav_burstcount -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata;                            // pixel_buffer_dma_0_avalon_pixel_dma_master_translator:uav_writedata -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_address;                              // pixel_buffer_dma_0_avalon_pixel_dma_master_translator:uav_address -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire          pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock;                                 // pixel_buffer_dma_0_avalon_pixel_dma_master_translator:uav_lock -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire          pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_write;                                // pixel_buffer_dma_0_avalon_pixel_dma_master_translator:uav_write -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire          pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_read;                                 // pixel_buffer_dma_0_avalon_pixel_dma_master_translator:uav_read -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata;                             // pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator:uav_readdata
	wire          pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess;                          // pixel_buffer_dma_0_avalon_pixel_dma_master_translator:uav_debugaccess -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable;                           // pixel_buffer_dma_0_avalon_pixel_dma_master_translator:uav_byteenable -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid;                        // pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator:uav_readdatavalid
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // nios2_processor_jtag_debug_module_translator:uav_waitrequest -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_processor_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                             // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_processor_jtag_debug_module_translator:uav_writedata
	wire   [31:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                               // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_processor_jtag_debug_module_translator:uav_address
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                 // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_processor_jtag_debug_module_translator:uav_write
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                  // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_processor_jtag_debug_module_translator:uav_lock
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                  // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_processor_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                              // nios2_processor_jtag_debug_module_translator:uav_readdata -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // nios2_processor_jtag_debug_module_translator:uav_readdatavalid -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_processor_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_processor_jtag_debug_module_translator:uav_byteenable
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                           // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                    // sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                     // sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                      // sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                        // sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                          // sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                           // sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                           // sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                       // sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                  // sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                    // sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                     // sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                             // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                   // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                           // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                    // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                   // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                          // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                        // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                 // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                // sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                              // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                               // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                              // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                                        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                    // timer_s1_translator:uav_waitrequest -> timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                     // timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_s1_translator:uav_burstcount
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                      // timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_s1_translator:uav_writedata
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                        // timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_s1_translator:uav_address
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                          // timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_s1_translator:uav_write
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                           // timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_s1_translator:uav_lock
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                           // timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_s1_translator:uav_read
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                       // timer_s1_translator:uav_readdata -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                  // timer_s1_translator:uav_readdatavalid -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                    // timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_s1_translator:uav_debugaccess
	wire    [3:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                     // timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_s1_translator:uav_byteenable
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                             // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                   // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                           // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                    // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                   // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                          // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                        // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                 // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                // timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                              // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                               // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                              // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // timestamp_s1_translator:uav_waitrequest -> timestamp_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timestamp_s1_translator:uav_burstcount
	wire   [31:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timestamp_s1_translator:uav_writedata
	wire   [31:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_address -> timestamp_s1_translator:uav_address
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_write -> timestamp_s1_translator:uav_write
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timestamp_s1_translator:uav_lock
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_read -> timestamp_s1_translator:uav_read
	wire   [31:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // timestamp_s1_translator:uav_readdata -> timestamp_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // timestamp_s1_translator:uav_readdatavalid -> timestamp_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timestamp_s1_translator:uav_debugaccess
	wire    [3:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timestamp_s1_translator:uav_byteenable
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // pixel_buffer_avalon_sram_slave_translator:uav_waitrequest -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> pixel_buffer_avalon_sram_slave_translator:uav_burstcount
	wire   [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> pixel_buffer_avalon_sram_slave_translator:uav_writedata
	wire   [31:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address;                                  // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> pixel_buffer_avalon_sram_slave_translator:uav_address
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write;                                    // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> pixel_buffer_avalon_sram_slave_translator:uav_write
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                     // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> pixel_buffer_avalon_sram_slave_translator:uav_lock
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read;                                     // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> pixel_buffer_avalon_sram_slave_translator:uav_read
	wire   [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // pixel_buffer_avalon_sram_slave_translator:uav_readdata -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // pixel_buffer_avalon_sram_slave_translator:uav_readdatavalid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pixel_buffer_avalon_sram_slave_translator:uav_debugaccess
	wire    [1:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> pixel_buffer_avalon_sram_slave_translator:uav_byteenable
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                              // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // pixel_buffer_dma_0_avalon_control_slave_translator:uav_waitrequest -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> pixel_buffer_dma_0_avalon_control_slave_translator:uav_burstcount
	wire   [31:0] pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                       // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> pixel_buffer_dma_0_avalon_control_slave_translator:uav_writedata
	wire   [31:0] pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                         // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> pixel_buffer_dma_0_avalon_control_slave_translator:uav_address
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                           // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> pixel_buffer_dma_0_avalon_control_slave_translator:uav_write
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                            // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> pixel_buffer_dma_0_avalon_control_slave_translator:uav_lock
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                            // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> pixel_buffer_dma_0_avalon_control_slave_translator:uav_read
	wire   [31:0] pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                        // pixel_buffer_dma_0_avalon_control_slave_translator:uav_readdata -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // pixel_buffer_dma_0_avalon_control_slave_translator:uav_readdatavalid -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pixel_buffer_dma_0_avalon_control_slave_translator:uav_debugaccess
	wire    [3:0] pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> pixel_buffer_dma_0_avalon_control_slave_translator:uav_byteenable
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                     // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // char_drawer_avalon_char_control_slave_translator:uav_waitrequest -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> char_drawer_avalon_char_control_slave_translator:uav_burstcount
	wire   [31:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                         // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> char_drawer_avalon_char_control_slave_translator:uav_writedata
	wire   [31:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                           // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> char_drawer_avalon_char_control_slave_translator:uav_address
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                             // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> char_drawer_avalon_char_control_slave_translator:uav_write
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                              // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> char_drawer_avalon_char_control_slave_translator:uav_lock
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                              // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> char_drawer_avalon_char_control_slave_translator:uav_read
	wire   [31:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                          // char_drawer_avalon_char_control_slave_translator:uav_readdata -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // char_drawer_avalon_char_control_slave_translator:uav_readdatavalid -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> char_drawer_avalon_char_control_slave_translator:uav_debugaccess
	wire    [3:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> char_drawer_avalon_char_control_slave_translator:uav_byteenable
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                       // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // char_drawer_avalon_char_buffer_slave_translator:uav_waitrequest -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> char_drawer_avalon_char_buffer_slave_translator:uav_burstcount
	wire    [7:0] char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> char_drawer_avalon_char_buffer_slave_translator:uav_writedata
	wire   [31:0] char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_address -> char_drawer_avalon_char_buffer_slave_translator:uav_address
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_write -> char_drawer_avalon_char_buffer_slave_translator:uav_write
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_lock -> char_drawer_avalon_char_buffer_slave_translator:uav_lock
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_read -> char_drawer_avalon_char_buffer_slave_translator:uav_read
	wire    [7:0] char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // char_drawer_avalon_char_buffer_slave_translator:uav_readdata -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // char_drawer_avalon_char_buffer_slave_translator:uav_readdatavalid -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> char_drawer_avalon_char_buffer_slave_translator:uav_debugaccess
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> char_drawer_avalon_char_buffer_slave_translator:uav_byteenable
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [80:0] char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [80:0] char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [7:0] char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                     // leds_s1_translator:uav_waitrequest -> leds_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                      // leds_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> leds_s1_translator:uav_burstcount
	wire   [31:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                       // leds_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> leds_s1_translator:uav_writedata
	wire   [31:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                         // leds_s1_translator_avalon_universal_slave_0_agent:m0_address -> leds_s1_translator:uav_address
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                           // leds_s1_translator_avalon_universal_slave_0_agent:m0_write -> leds_s1_translator:uav_write
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                            // leds_s1_translator_avalon_universal_slave_0_agent:m0_lock -> leds_s1_translator:uav_lock
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                            // leds_s1_translator_avalon_universal_slave_0_agent:m0_read -> leds_s1_translator:uav_read
	wire   [31:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                        // leds_s1_translator:uav_readdata -> leds_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                   // leds_s1_translator:uav_readdatavalid -> leds_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                     // leds_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> leds_s1_translator:uav_debugaccess
	wire    [3:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                      // leds_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> leds_s1_translator:uav_byteenable
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                              // leds_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                    // leds_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                            // leds_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                     // leds_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                    // leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> leds_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                           // leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                 // leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                         // leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                  // leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                 // leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                               // leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                // leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                               // leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // SD_Card_avalon_sdcard_slave_translator:uav_waitrequest -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> SD_Card_avalon_sdcard_slave_translator:uav_burstcount
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> SD_Card_avalon_sdcard_slave_translator:uav_writedata
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address;                                     // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_address -> SD_Card_avalon_sdcard_slave_translator:uav_address
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write;                                       // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_write -> SD_Card_avalon_sdcard_slave_translator:uav_write
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                        // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_lock -> SD_Card_avalon_sdcard_slave_translator:uav_lock
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read;                                        // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_read -> SD_Card_avalon_sdcard_slave_translator:uav_read
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // SD_Card_avalon_sdcard_slave_translator:uav_readdata -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // SD_Card_avalon_sdcard_slave_translator:uav_readdatavalid -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SD_Card_avalon_sdcard_slave_translator:uav_debugaccess
	wire    [3:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> SD_Card_avalon_sdcard_slave_translator:uav_byteenable
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                 // Switches_s1_translator:uav_waitrequest -> Switches_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                  // Switches_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> Switches_s1_translator:uav_burstcount
	wire   [31:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                   // Switches_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> Switches_s1_translator:uav_writedata
	wire   [31:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                     // Switches_s1_translator_avalon_universal_slave_0_agent:m0_address -> Switches_s1_translator:uav_address
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                       // Switches_s1_translator_avalon_universal_slave_0_agent:m0_write -> Switches_s1_translator:uav_write
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                        // Switches_s1_translator_avalon_universal_slave_0_agent:m0_lock -> Switches_s1_translator:uav_lock
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                        // Switches_s1_translator_avalon_universal_slave_0_agent:m0_read -> Switches_s1_translator:uav_read
	wire   [31:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                    // Switches_s1_translator:uav_readdata -> Switches_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                               // Switches_s1_translator:uav_readdatavalid -> Switches_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                 // Switches_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Switches_s1_translator:uav_debugaccess
	wire    [3:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                  // Switches_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> Switches_s1_translator:uav_byteenable
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                          // Switches_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                // Switches_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                        // Switches_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] switches_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                 // Switches_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                // Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Switches_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                       // Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                             // Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                     // Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                              // Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                             // Switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                           // Switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                            // Switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                           // Switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          keys_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                     // Keys_s1_translator:uav_waitrequest -> Keys_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] keys_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                      // Keys_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> Keys_s1_translator:uav_burstcount
	wire   [31:0] keys_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                       // Keys_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> Keys_s1_translator:uav_writedata
	wire   [31:0] keys_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                         // Keys_s1_translator_avalon_universal_slave_0_agent:m0_address -> Keys_s1_translator:uav_address
	wire          keys_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                           // Keys_s1_translator_avalon_universal_slave_0_agent:m0_write -> Keys_s1_translator:uav_write
	wire          keys_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                            // Keys_s1_translator_avalon_universal_slave_0_agent:m0_lock -> Keys_s1_translator:uav_lock
	wire          keys_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                            // Keys_s1_translator_avalon_universal_slave_0_agent:m0_read -> Keys_s1_translator:uav_read
	wire   [31:0] keys_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                        // Keys_s1_translator:uav_readdata -> Keys_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          keys_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                   // Keys_s1_translator:uav_readdatavalid -> Keys_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          keys_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                     // Keys_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Keys_s1_translator:uav_debugaccess
	wire    [3:0] keys_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                      // Keys_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> Keys_s1_translator:uav_byteenable
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                              // Keys_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                    // Keys_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> Keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                            // Keys_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] keys_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                     // Keys_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> Keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                    // Keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Keys_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                           // Keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Keys_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                 // Keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Keys_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                         // Keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Keys_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                  // Keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Keys_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                 // Keys_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                               // Keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                // Keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                               // Keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // audio_and_video_config_0_avalon_av_config_slave_translator:uav_waitrequest -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_burstcount
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_writedata
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_address -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_address
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_write -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_write
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_lock -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_lock
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_read -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_read
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // audio_and_video_config_0_avalon_av_config_slave_translator:uav_readdata -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // audio_and_video_config_0_avalon_av_config_slave_translator:uav_readdatavalid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_debugaccess
	wire    [3:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_byteenable
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // audio_avalon_audio_slave_translator:uav_waitrequest -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_avalon_audio_slave_translator:uav_burstcount
	wire   [31:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_avalon_audio_slave_translator:uav_writedata
	wire   [31:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_address;                                        // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_address -> audio_avalon_audio_slave_translator:uav_address
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_write;                                          // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_write -> audio_avalon_audio_slave_translator:uav_write
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                           // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_lock -> audio_avalon_audio_slave_translator:uav_lock
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_read;                                           // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_read -> audio_avalon_audio_slave_translator:uav_read
	wire   [31:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // audio_avalon_audio_slave_translator:uav_readdata -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // audio_avalon_audio_slave_translator:uav_readdatavalid -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_avalon_audio_slave_translator:uav_debugaccess
	wire    [3:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_avalon_audio_slave_translator:uav_byteenable
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                     // LEDR_s1_translator:uav_waitrequest -> LEDR_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                      // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LEDR_s1_translator:uav_burstcount
	wire   [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                       // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LEDR_s1_translator:uav_writedata
	wire   [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                         // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_address -> LEDR_s1_translator:uav_address
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                           // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_write -> LEDR_s1_translator:uav_write
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                            // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LEDR_s1_translator:uav_lock
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                            // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_read -> LEDR_s1_translator:uav_read
	wire   [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                        // LEDR_s1_translator:uav_readdata -> LEDR_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                   // LEDR_s1_translator:uav_readdatavalid -> LEDR_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                     // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LEDR_s1_translator:uav_debugaccess
	wire    [3:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                      // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LEDR_s1_translator:uav_byteenable
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                              // LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                    // LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                            // LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                     // LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                    // LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                           // LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                 // LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                         // LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                  // LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                 // LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                               // LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                // LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                               // LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // ps2_0_avalon_ps2_slave_translator:uav_waitrequest -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> ps2_0_avalon_ps2_slave_translator:uav_burstcount
	wire   [31:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> ps2_0_avalon_ps2_slave_translator:uav_writedata
	wire   [31:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_address;                                          // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_address -> ps2_0_avalon_ps2_slave_translator:uav_address
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_write;                                            // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_write -> ps2_0_avalon_ps2_slave_translator:uav_write
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                             // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_lock -> ps2_0_avalon_ps2_slave_translator:uav_lock
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_read;                                             // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_read -> ps2_0_avalon_ps2_slave_translator:uav_read
	wire   [31:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // ps2_0_avalon_ps2_slave_translator:uav_readdata -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // ps2_0_avalon_ps2_slave_translator:uav_readdatavalid -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ps2_0_avalon_ps2_slave_translator:uav_debugaccess
	wire    [3:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> ps2_0_avalon_ps2_slave_translator:uav_byteenable
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                     // hex0_s1_translator:uav_waitrequest -> hex0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hex0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                      // hex0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex0_s1_translator:uav_burstcount
	wire   [31:0] hex0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                       // hex0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex0_s1_translator:uav_writedata
	wire   [31:0] hex0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                         // hex0_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex0_s1_translator:uav_address
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                           // hex0_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex0_s1_translator:uav_write
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                            // hex0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex0_s1_translator:uav_lock
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                            // hex0_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex0_s1_translator:uav_read
	wire   [31:0] hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                        // hex0_s1_translator:uav_readdata -> hex0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                   // hex0_s1_translator:uav_readdatavalid -> hex0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                     // hex0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex0_s1_translator:uav_debugaccess
	wire    [3:0] hex0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                      // hex0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex0_s1_translator:uav_byteenable
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                              // hex0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                    // hex0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                            // hex0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                     // hex0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                    // hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                           // hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                 // hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                         // hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                  // hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                 // hex0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                               // hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                // hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                               // hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                     // hex1_s1_translator:uav_waitrequest -> hex1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hex1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                      // hex1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex1_s1_translator:uav_burstcount
	wire   [31:0] hex1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                       // hex1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex1_s1_translator:uav_writedata
	wire   [31:0] hex1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                         // hex1_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex1_s1_translator:uav_address
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                           // hex1_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex1_s1_translator:uav_write
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                            // hex1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex1_s1_translator:uav_lock
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                            // hex1_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex1_s1_translator:uav_read
	wire   [31:0] hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                        // hex1_s1_translator:uav_readdata -> hex1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                   // hex1_s1_translator:uav_readdatavalid -> hex1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                     // hex1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex1_s1_translator:uav_debugaccess
	wire    [3:0] hex1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                      // hex1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex1_s1_translator:uav_byteenable
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                              // hex1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                    // hex1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                            // hex1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                     // hex1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                    // hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                           // hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                 // hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                         // hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                  // hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                 // hex1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                               // hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                // hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                               // hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                     // hex2_s1_translator:uav_waitrequest -> hex2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hex2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                      // hex2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex2_s1_translator:uav_burstcount
	wire   [31:0] hex2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                       // hex2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex2_s1_translator:uav_writedata
	wire   [31:0] hex2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                         // hex2_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex2_s1_translator:uav_address
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                           // hex2_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex2_s1_translator:uav_write
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                            // hex2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex2_s1_translator:uav_lock
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                            // hex2_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex2_s1_translator:uav_read
	wire   [31:0] hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                        // hex2_s1_translator:uav_readdata -> hex2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                   // hex2_s1_translator:uav_readdatavalid -> hex2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                     // hex2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex2_s1_translator:uav_debugaccess
	wire    [3:0] hex2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                      // hex2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex2_s1_translator:uav_byteenable
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                              // hex2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                    // hex2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                            // hex2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                     // hex2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                    // hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                           // hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                 // hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                         // hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                  // hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                 // hex2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                               // hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                // hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                               // hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                     // hex3_s1_translator:uav_waitrequest -> hex3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hex3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                      // hex3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex3_s1_translator:uav_burstcount
	wire   [31:0] hex3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                       // hex3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex3_s1_translator:uav_writedata
	wire   [31:0] hex3_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                         // hex3_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex3_s1_translator:uav_address
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                           // hex3_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex3_s1_translator:uav_write
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                            // hex3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex3_s1_translator:uav_lock
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                            // hex3_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex3_s1_translator:uav_read
	wire   [31:0] hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                        // hex3_s1_translator:uav_readdata -> hex3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                   // hex3_s1_translator:uav_readdatavalid -> hex3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                     // hex3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex3_s1_translator:uav_debugaccess
	wire    [3:0] hex3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                      // hex3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex3_s1_translator:uav_byteenable
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                              // hex3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                    // hex3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                            // hex3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                     // hex3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                    // hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                           // hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                 // hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                         // hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                  // hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                 // hex3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                               // hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                // hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                               // hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                     // hex4_s1_translator:uav_waitrequest -> hex4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hex4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                      // hex4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex4_s1_translator:uav_burstcount
	wire   [31:0] hex4_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                       // hex4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex4_s1_translator:uav_writedata
	wire   [31:0] hex4_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                         // hex4_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex4_s1_translator:uav_address
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                           // hex4_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex4_s1_translator:uav_write
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                            // hex4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex4_s1_translator:uav_lock
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                            // hex4_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex4_s1_translator:uav_read
	wire   [31:0] hex4_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                        // hex4_s1_translator:uav_readdata -> hex4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                   // hex4_s1_translator:uav_readdatavalid -> hex4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                     // hex4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex4_s1_translator:uav_debugaccess
	wire    [3:0] hex4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                      // hex4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex4_s1_translator:uav_byteenable
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                              // hex4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                    // hex4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                            // hex4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                     // hex4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                    // hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                           // hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                 // hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                         // hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                  // hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                 // hex4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                               // hex4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                // hex4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                               // hex4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // character_lcd_0_avalon_lcd_slave_translator:uav_waitrequest -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> character_lcd_0_avalon_lcd_slave_translator:uav_burstcount
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                              // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> character_lcd_0_avalon_lcd_slave_translator:uav_writedata
	wire   [31:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address;                                // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_address -> character_lcd_0_avalon_lcd_slave_translator:uav_address
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write;                                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_write -> character_lcd_0_avalon_lcd_slave_translator:uav_write
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                   // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_lock -> character_lcd_0_avalon_lcd_slave_translator:uav_lock
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read;                                   // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_read -> character_lcd_0_avalon_lcd_slave_translator:uav_read
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                               // character_lcd_0_avalon_lcd_slave_translator:uav_readdata -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // character_lcd_0_avalon_lcd_slave_translator:uav_readdatavalid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> character_lcd_0_avalon_lcd_slave_translator:uav_debugaccess
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> character_lcd_0_avalon_lcd_slave_translator:uav_byteenable
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [80:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [80:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                         // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                               // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                       // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [106:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                                // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                               // addr_router:sink_ready -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                // nios2_processor_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                      // nios2_processor_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                              // nios2_processor_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [106:0] nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_data;                                       // nios2_processor_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                      // addr_router_001:sink_ready -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid;                       // pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire   [88:0] pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data;                        // pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_002:sink_ready -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                 // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [106:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                  // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router:sink_ready -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                    // sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                          // sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                  // sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [88:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                           // sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                          // id_router_001:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [106:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                                        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_002:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                    // timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                          // timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                  // timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [106:0] timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                           // timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                          // id_router_003:sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [106:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_004:sink_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                    // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire   [88:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data;                                     // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_005:sink_ready -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                           // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [106:0] pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                            // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_006:sink_ready -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                             // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [106:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                              // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_007:sink_ready -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire   [79:0] char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_008:sink_ready -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                     // leds_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                           // leds_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                   // leds_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [106:0] leds_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                            // leds_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                           // id_router_009:sink_ready -> leds_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                       // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [106:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data;                                        // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_010:sink_ready -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                 // Switches_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                       // Switches_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                               // Switches_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [106:0] switches_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                        // Switches_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                       // id_router_011:sink_ready -> Switches_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                     // Keys_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                           // Keys_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                   // Keys_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [106:0] keys_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                            // Keys_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                           // id_router_012:sink_ready -> Keys_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [106:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_013:sink_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                          // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [106:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_data;                                           // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_014:sink_ready -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                     // LEDR_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                           // LEDR_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                   // LEDR_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [106:0] ledr_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                            // LEDR_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                           // id_router_015:sink_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                            // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [106:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_data;                                             // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_016:sink_ready -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                     // hex0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                           // hex0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                   // hex0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [106:0] hex0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                            // hex0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                           // id_router_017:sink_ready -> hex0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                     // hex1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                           // hex1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                   // hex1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [106:0] hex1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                            // hex1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                           // id_router_018:sink_ready -> hex1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                     // hex2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                           // hex2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                   // hex2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire  [106:0] hex2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                            // hex2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                           // id_router_019:sink_ready -> hex2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                     // hex3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                           // hex3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                   // hex3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire  [106:0] hex3_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                            // hex3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                           // id_router_020:sink_ready -> hex3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                     // hex4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                           // hex4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                   // hex4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire  [106:0] hex4_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                            // hex4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire          hex4_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                           // id_router_021:sink_ready -> hex4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	wire   [79:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data;                                   // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_022:sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                                          // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                                                // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                                        // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [106:0] addr_router_src_data;                                                                                                 // addr_router:src_data -> limiter:cmd_sink_data
	wire   [22:0] addr_router_src_channel;                                                                                              // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                                                // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                                          // limiter:rsp_src_endofpacket -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                                // limiter:rsp_src_valid -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                                        // limiter:rsp_src_startofpacket -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_rsp_src_data;                                                                                                 // limiter:rsp_src_data -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [22:0] limiter_rsp_src_channel;                                                                                              // limiter:rsp_src_channel -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                                // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_001_src_endofpacket;                                                                                      // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                            // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_001_src_startofpacket;                                                                                    // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [106:0] addr_router_001_src_data;                                                                                             // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire   [22:0] addr_router_001_src_channel;                                                                                          // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_001_src_ready;                                                                                            // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                                      // limiter_001:rsp_src_endofpacket -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                                            // limiter_001:rsp_src_valid -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                                    // limiter_001:rsp_src_startofpacket -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_001_rsp_src_data;                                                                                             // limiter_001:rsp_src_data -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [22:0] limiter_001_rsp_src_channel;                                                                                          // limiter_001:rsp_src_channel -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                                            // nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                                    // burst_adapter:source0_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                                          // burst_adapter:source0_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                                  // burst_adapter:source0_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] burst_adapter_source0_data;                                                                                           // burst_adapter:source0_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                                          // sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [22:0] burst_adapter_source0_channel;                                                                                        // burst_adapter:source0_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                                                // burst_adapter_001:source0_endofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                                      // burst_adapter_001:source0_valid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                                              // burst_adapter_001:source0_startofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] burst_adapter_001_source0_data;                                                                                       // burst_adapter_001:source0_data -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                                      // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [22:0] burst_adapter_001_source0_channel;                                                                                    // burst_adapter_001:source0_channel -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_002_source0_endofpacket;                                                                                // burst_adapter_002:source0_endofpacket -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_002_source0_valid;                                                                                      // burst_adapter_002:source0_valid -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_002_source0_startofpacket;                                                                              // burst_adapter_002:source0_startofpacket -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [79:0] burst_adapter_002_source0_data;                                                                                       // burst_adapter_002:source0_data -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_002_source0_ready;                                                                                      // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire   [22:0] burst_adapter_002_source0_channel;                                                                                    // burst_adapter_002:source0_channel -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_003_source0_endofpacket;                                                                                // burst_adapter_003:source0_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_003_source0_valid;                                                                                      // burst_adapter_003:source0_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_003_source0_startofpacket;                                                                              // burst_adapter_003:source0_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [79:0] burst_adapter_003_source0_data;                                                                                       // burst_adapter_003:source0_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_003_source0_ready;                                                                                      // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	wire   [22:0] burst_adapter_003_source0_channel;                                                                                    // burst_adapter_003:source0_channel -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                                       // rst_controller:reset_out -> [Keys:reset_n, Keys_s1_translator:reset, Keys_s1_translator_avalon_universal_slave_0_agent:reset, Keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LEDR:reset_n, LEDR_s1_translator:reset, LEDR_s1_translator_avalon_universal_slave_0_agent:reset, LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SD_Card:i_reset_n, SD_Card_avalon_sdcard_slave_translator:reset, SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:reset, SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Switches:reset_n, Switches_s1_translator:reset, Switches_s1_translator_avalon_universal_slave_0_agent:reset, Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, addr_router_002:reset, alpha_blender:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, burst_adapter_003:reset, char_drawer:reset, char_drawer_avalon_char_buffer_slave_translator:reset, char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:reset, char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, char_drawer_avalon_char_control_slave_translator:reset, char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:reset, char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, character_lcd_0:reset, character_lcd_0_avalon_lcd_slave_translator:reset, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:reset, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_005:reset, hex0:reset_n, hex0_s1_translator:reset, hex0_s1_translator_avalon_universal_slave_0_agent:reset, hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hex1:reset_n, hex1_s1_translator:reset, hex1_s1_translator_avalon_universal_slave_0_agent:reset, hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hex2:reset_n, hex2_s1_translator:reset, hex2_s1_translator_avalon_universal_slave_0_agent:reset, hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hex3:reset_n, hex3_s1_translator:reset, hex3_s1_translator_avalon_universal_slave_0_agent:reset, hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hex4:reset_n, hex4_s1_translator:reset, hex4_s1_translator_avalon_universal_slave_0_agent:reset, hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, id_router_022:reset, irq_mapper:reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, leds:reset_n, leds_s1_translator:reset, leds_s1_translator_avalon_universal_slave_0_agent:reset, leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, nios2_processor:reset_n, nios2_processor_data_master_translator:reset, nios2_processor_data_master_translator_avalon_universal_master_0_agent:reset, nios2_processor_instruction_master_translator:reset, nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_processor_jtag_debug_module_translator:reset, nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pixel_buffer:reset, pixel_buffer_avalon_sram_slave_translator:reset, pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pixel_buffer_dma_0:reset, pixel_buffer_dma_0_avalon_control_slave_translator:reset, pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:reset, pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pixel_buffer_dma_0_avalon_pixel_dma_master_translator:reset, pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:reset, ps2_0:reset, ps2_0_avalon_ps2_slave_translator:reset, ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:reset, ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rgb_resampler:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_022:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, scaler:reset, sdram:reset_n, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer:reset_n, timer_s1_translator:reset, timer_s1_translator_avalon_universal_slave_0_agent:reset, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timestamp:reset_n, timestamp_s1_translator:reset, timestamp_s1_translator_avalon_universal_slave_0_agent:reset, timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, video_fifo:reset_stream_in, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset, width_adapter_008:reset, width_adapter_009:reset]
	wire          nios2_processor_jtag_debug_module_reset_reset;                                                                        // nios2_processor:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	wire          rst_controller_001_reset_out_reset;                                                                                   // rst_controller_001:reset_out -> clocks:reset
	wire          rst_controller_002_reset_out_reset;                                                                                   // rst_controller_002:reset_out -> [vga_controller:reset, video_fifo:reset_stream_out]
	wire          rst_controller_003_reset_out_reset;                                                                                   // rst_controller_003:reset_out -> [audio:reset, audio_and_video_config_0:reset, audio_and_video_config_0_avalon_av_config_slave_translator:reset, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:reset, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, audio_avalon_audio_slave_translator:reset, audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:reset, audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_013:reset, id_router_014:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, up_clocks_0:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                                      // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                            // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                                    // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src0_data;                                                                                             // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [22:0] cmd_xbar_demux_src0_channel;                                                                                          // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                            // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                                  // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                                        // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                                // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src0_data;                                                                                         // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [22:0] cmd_xbar_demux_001_src0_channel;                                                                                      // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                                        // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                                  // cmd_xbar_demux_001:src2_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                                        // cmd_xbar_demux_001:src2_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                                // cmd_xbar_demux_001:src2_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src2_data;                                                                                         // cmd_xbar_demux_001:src2_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src2_channel;                                                                                      // cmd_xbar_demux_001:src2_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                                  // cmd_xbar_demux_001:src3_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                                        // cmd_xbar_demux_001:src3_valid -> timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                                // cmd_xbar_demux_001:src3_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src3_data;                                                                                         // cmd_xbar_demux_001:src3_data -> timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src3_channel;                                                                                      // cmd_xbar_demux_001:src3_channel -> timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                                  // cmd_xbar_demux_001:src4_endofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                                        // cmd_xbar_demux_001:src4_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                                // cmd_xbar_demux_001:src4_startofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src4_data;                                                                                         // cmd_xbar_demux_001:src4_data -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src4_channel;                                                                                      // cmd_xbar_demux_001:src4_channel -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                                  // cmd_xbar_demux_001:src6_endofpacket -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                                        // cmd_xbar_demux_001:src6_valid -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                                // cmd_xbar_demux_001:src6_startofpacket -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src6_data;                                                                                         // cmd_xbar_demux_001:src6_data -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src6_channel;                                                                                      // cmd_xbar_demux_001:src6_channel -> pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                                  // cmd_xbar_demux_001:src7_endofpacket -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                                        // cmd_xbar_demux_001:src7_valid -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                                // cmd_xbar_demux_001:src7_startofpacket -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src7_data;                                                                                         // cmd_xbar_demux_001:src7_data -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src7_channel;                                                                                      // cmd_xbar_demux_001:src7_channel -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                                                  // cmd_xbar_demux_001:src9_endofpacket -> leds_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                                        // cmd_xbar_demux_001:src9_valid -> leds_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                                                // cmd_xbar_demux_001:src9_startofpacket -> leds_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src9_data;                                                                                         // cmd_xbar_demux_001:src9_data -> leds_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src9_channel;                                                                                      // cmd_xbar_demux_001:src9_channel -> leds_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                                                 // cmd_xbar_demux_001:src10_endofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                                       // cmd_xbar_demux_001:src10_valid -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                                               // cmd_xbar_demux_001:src10_startofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src10_data;                                                                                        // cmd_xbar_demux_001:src10_data -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src10_channel;                                                                                     // cmd_xbar_demux_001:src10_channel -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                                                 // cmd_xbar_demux_001:src11_endofpacket -> Switches_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                                       // cmd_xbar_demux_001:src11_valid -> Switches_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                                               // cmd_xbar_demux_001:src11_startofpacket -> Switches_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src11_data;                                                                                        // cmd_xbar_demux_001:src11_data -> Switches_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src11_channel;                                                                                     // cmd_xbar_demux_001:src11_channel -> Switches_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src12_endofpacket;                                                                                 // cmd_xbar_demux_001:src12_endofpacket -> Keys_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src12_valid;                                                                                       // cmd_xbar_demux_001:src12_valid -> Keys_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src12_startofpacket;                                                                               // cmd_xbar_demux_001:src12_startofpacket -> Keys_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src12_data;                                                                                        // cmd_xbar_demux_001:src12_data -> Keys_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src12_channel;                                                                                     // cmd_xbar_demux_001:src12_channel -> Keys_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src13_endofpacket;                                                                                 // cmd_xbar_demux_001:src13_endofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src13_valid;                                                                                       // cmd_xbar_demux_001:src13_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src13_startofpacket;                                                                               // cmd_xbar_demux_001:src13_startofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src13_data;                                                                                        // cmd_xbar_demux_001:src13_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src13_channel;                                                                                     // cmd_xbar_demux_001:src13_channel -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src14_endofpacket;                                                                                 // cmd_xbar_demux_001:src14_endofpacket -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src14_valid;                                                                                       // cmd_xbar_demux_001:src14_valid -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src14_startofpacket;                                                                               // cmd_xbar_demux_001:src14_startofpacket -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src14_data;                                                                                        // cmd_xbar_demux_001:src14_data -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src14_channel;                                                                                     // cmd_xbar_demux_001:src14_channel -> audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src15_endofpacket;                                                                                 // cmd_xbar_demux_001:src15_endofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src15_valid;                                                                                       // cmd_xbar_demux_001:src15_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src15_startofpacket;                                                                               // cmd_xbar_demux_001:src15_startofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src15_data;                                                                                        // cmd_xbar_demux_001:src15_data -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src15_channel;                                                                                     // cmd_xbar_demux_001:src15_channel -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src16_endofpacket;                                                                                 // cmd_xbar_demux_001:src16_endofpacket -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src16_valid;                                                                                       // cmd_xbar_demux_001:src16_valid -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src16_startofpacket;                                                                               // cmd_xbar_demux_001:src16_startofpacket -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src16_data;                                                                                        // cmd_xbar_demux_001:src16_data -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src16_channel;                                                                                     // cmd_xbar_demux_001:src16_channel -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src17_endofpacket;                                                                                 // cmd_xbar_demux_001:src17_endofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src17_valid;                                                                                       // cmd_xbar_demux_001:src17_valid -> hex0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src17_startofpacket;                                                                               // cmd_xbar_demux_001:src17_startofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src17_data;                                                                                        // cmd_xbar_demux_001:src17_data -> hex0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src17_channel;                                                                                     // cmd_xbar_demux_001:src17_channel -> hex0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src18_endofpacket;                                                                                 // cmd_xbar_demux_001:src18_endofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src18_valid;                                                                                       // cmd_xbar_demux_001:src18_valid -> hex1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src18_startofpacket;                                                                               // cmd_xbar_demux_001:src18_startofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src18_data;                                                                                        // cmd_xbar_demux_001:src18_data -> hex1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src18_channel;                                                                                     // cmd_xbar_demux_001:src18_channel -> hex1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src19_endofpacket;                                                                                 // cmd_xbar_demux_001:src19_endofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src19_valid;                                                                                       // cmd_xbar_demux_001:src19_valid -> hex2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src19_startofpacket;                                                                               // cmd_xbar_demux_001:src19_startofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src19_data;                                                                                        // cmd_xbar_demux_001:src19_data -> hex2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src19_channel;                                                                                     // cmd_xbar_demux_001:src19_channel -> hex2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src20_endofpacket;                                                                                 // cmd_xbar_demux_001:src20_endofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src20_valid;                                                                                       // cmd_xbar_demux_001:src20_valid -> hex3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src20_startofpacket;                                                                               // cmd_xbar_demux_001:src20_startofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src20_data;                                                                                        // cmd_xbar_demux_001:src20_data -> hex3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src20_channel;                                                                                     // cmd_xbar_demux_001:src20_channel -> hex3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src21_endofpacket;                                                                                 // cmd_xbar_demux_001:src21_endofpacket -> hex4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src21_valid;                                                                                       // cmd_xbar_demux_001:src21_valid -> hex4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src21_startofpacket;                                                                               // cmd_xbar_demux_001:src21_startofpacket -> hex4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src21_data;                                                                                        // cmd_xbar_demux_001:src21_data -> hex4_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src21_channel;                                                                                     // cmd_xbar_demux_001:src21_channel -> hex4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                                  // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                                        // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_005:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                                // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire   [88:0] cmd_xbar_demux_002_src0_data;                                                                                         // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_005:sink1_data
	wire   [22:0] cmd_xbar_demux_002_src0_channel;                                                                                      // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_005:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                                        // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                                      // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                            // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                                    // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_src0_data;                                                                                             // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [22:0] rsp_xbar_demux_src0_channel;                                                                                          // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                            // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                                      // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                            // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                                    // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_src1_data;                                                                                             // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [22:0] rsp_xbar_demux_src1_channel;                                                                                          // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                            // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                                  // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                                        // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                                // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_002_src0_data;                                                                                         // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	wire   [22:0] rsp_xbar_demux_002_src0_channel;                                                                                      // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                                        // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                                  // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                                        // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                                // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src0_data;                                                                                         // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [22:0] rsp_xbar_demux_003_src0_channel;                                                                                      // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                                        // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                                  // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                                        // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                                // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [106:0] rsp_xbar_demux_004_src0_data;                                                                                         // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [22:0] rsp_xbar_demux_004_src0_channel;                                                                                      // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                                        // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src1_endofpacket;                                                                                  // rsp_xbar_demux_005:src1_endofpacket -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_005_src1_valid;                                                                                        // rsp_xbar_demux_005:src1_valid -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_005_src1_startofpacket;                                                                                // rsp_xbar_demux_005:src1_startofpacket -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] rsp_xbar_demux_005_src1_data;                                                                                         // rsp_xbar_demux_005:src1_data -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [22:0] rsp_xbar_demux_005_src1_channel;                                                                                      // rsp_xbar_demux_005:src1_channel -> pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                                  // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                                        // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                                // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [106:0] rsp_xbar_demux_006_src0_data;                                                                                         // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [22:0] rsp_xbar_demux_006_src0_channel;                                                                                      // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                                        // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                                  // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                                        // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                                // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [106:0] rsp_xbar_demux_007_src0_data;                                                                                         // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [22:0] rsp_xbar_demux_007_src0_channel;                                                                                      // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                                        // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                                  // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                                        // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                                // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [106:0] rsp_xbar_demux_009_src0_data;                                                                                         // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire   [22:0] rsp_xbar_demux_009_src0_channel;                                                                                      // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                                        // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                                  // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                                        // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                                // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [106:0] rsp_xbar_demux_010_src0_data;                                                                                         // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire   [22:0] rsp_xbar_demux_010_src0_channel;                                                                                      // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                                        // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                                  // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                                        // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                                // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [106:0] rsp_xbar_demux_011_src0_data;                                                                                         // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire   [22:0] rsp_xbar_demux_011_src0_channel;                                                                                      // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                                        // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                                  // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                                        // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                                // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [106:0] rsp_xbar_demux_012_src0_data;                                                                                         // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire   [22:0] rsp_xbar_demux_012_src0_channel;                                                                                      // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                                        // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                                  // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                                        // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                                // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [106:0] rsp_xbar_demux_013_src0_data;                                                                                         // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	wire   [22:0] rsp_xbar_demux_013_src0_channel;                                                                                      // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                                        // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                                  // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                                        // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                                // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [106:0] rsp_xbar_demux_014_src0_data;                                                                                         // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	wire   [22:0] rsp_xbar_demux_014_src0_channel;                                                                                      // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                                        // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                                  // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                                        // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                                // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [106:0] rsp_xbar_demux_015_src0_data;                                                                                         // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	wire   [22:0] rsp_xbar_demux_015_src0_channel;                                                                                      // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                                        // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                                                  // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                                        // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_001:sink16_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                                                // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [106:0] rsp_xbar_demux_016_src0_data;                                                                                         // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_001:sink16_data
	wire   [22:0] rsp_xbar_demux_016_src0_channel;                                                                                      // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_001:sink16_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                                        // rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                                                  // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                                        // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_001:sink17_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                                                // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	wire  [106:0] rsp_xbar_demux_017_src0_data;                                                                                         // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_001:sink17_data
	wire   [22:0] rsp_xbar_demux_017_src0_channel;                                                                                      // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_001:sink17_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                                        // rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                                                  // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                                        // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_001:sink18_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                                                // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	wire  [106:0] rsp_xbar_demux_018_src0_data;                                                                                         // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_001:sink18_data
	wire   [22:0] rsp_xbar_demux_018_src0_channel;                                                                                      // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_001:sink18_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                                        // rsp_xbar_mux_001:sink18_ready -> rsp_xbar_demux_018:src0_ready
	wire          rsp_xbar_demux_019_src0_endofpacket;                                                                                  // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_001:sink19_endofpacket
	wire          rsp_xbar_demux_019_src0_valid;                                                                                        // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_001:sink19_valid
	wire          rsp_xbar_demux_019_src0_startofpacket;                                                                                // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_001:sink19_startofpacket
	wire  [106:0] rsp_xbar_demux_019_src0_data;                                                                                         // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_001:sink19_data
	wire   [22:0] rsp_xbar_demux_019_src0_channel;                                                                                      // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_001:sink19_channel
	wire          rsp_xbar_demux_019_src0_ready;                                                                                        // rsp_xbar_mux_001:sink19_ready -> rsp_xbar_demux_019:src0_ready
	wire          rsp_xbar_demux_020_src0_endofpacket;                                                                                  // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_001:sink20_endofpacket
	wire          rsp_xbar_demux_020_src0_valid;                                                                                        // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_001:sink20_valid
	wire          rsp_xbar_demux_020_src0_startofpacket;                                                                                // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_001:sink20_startofpacket
	wire  [106:0] rsp_xbar_demux_020_src0_data;                                                                                         // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_001:sink20_data
	wire   [22:0] rsp_xbar_demux_020_src0_channel;                                                                                      // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_001:sink20_channel
	wire          rsp_xbar_demux_020_src0_ready;                                                                                        // rsp_xbar_mux_001:sink20_ready -> rsp_xbar_demux_020:src0_ready
	wire          rsp_xbar_demux_021_src0_endofpacket;                                                                                  // rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_001:sink21_endofpacket
	wire          rsp_xbar_demux_021_src0_valid;                                                                                        // rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_001:sink21_valid
	wire          rsp_xbar_demux_021_src0_startofpacket;                                                                                // rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_001:sink21_startofpacket
	wire  [106:0] rsp_xbar_demux_021_src0_data;                                                                                         // rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_001:sink21_data
	wire   [22:0] rsp_xbar_demux_021_src0_channel;                                                                                      // rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_001:sink21_channel
	wire          rsp_xbar_demux_021_src0_ready;                                                                                        // rsp_xbar_mux_001:sink21_ready -> rsp_xbar_demux_021:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                                          // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                                        // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [106:0] limiter_cmd_src_data;                                                                                                 // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [22:0] limiter_cmd_src_channel;                                                                                              // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                                                // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                                         // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                               // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                                       // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_src_data;                                                                                                // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [22:0] rsp_xbar_mux_src_channel;                                                                                             // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                                               // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                                      // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                                    // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [106:0] limiter_001_cmd_src_data;                                                                                             // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire   [22:0] limiter_001_cmd_src_channel;                                                                                          // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                                            // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                                     // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                           // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                                   // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_001_src_data;                                                                                            // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire   [22:0] rsp_xbar_mux_001_src_channel;                                                                                         // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                           // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire          addr_router_002_src_endofpacket;                                                                                      // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                                            // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                                    // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire   [88:0] addr_router_002_src_data;                                                                                             // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire   [22:0] addr_router_002_src_channel;                                                                                          // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                                            // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_demux_005_src1_ready;                                                                                        // pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_005:src1_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                                         // cmd_xbar_mux:src_endofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                               // cmd_xbar_mux:src_valid -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                                       // cmd_xbar_mux:src_startofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_src_data;                                                                                                // cmd_xbar_mux:src_data -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_mux_src_channel;                                                                                             // cmd_xbar_mux:src_channel -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                               // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                            // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                                  // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                                          // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [106:0] id_router_src_data;                                                                                                   // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [22:0] id_router_src_channel;                                                                                                // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                                  // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                                     // cmd_xbar_mux_001:src_endofpacket -> burst_adapter:sink0_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                                           // cmd_xbar_mux_001:src_valid -> burst_adapter:sink0_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                                   // cmd_xbar_mux_001:src_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [88:0] cmd_xbar_mux_001_src_data;                                                                                            // cmd_xbar_mux_001:src_data -> burst_adapter:sink0_data
	wire   [22:0] cmd_xbar_mux_001_src_channel;                                                                                         // cmd_xbar_mux_001:src_channel -> burst_adapter:sink0_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                                           // burst_adapter:sink0_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                                        // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                              // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                                      // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire   [88:0] id_router_001_src_data;                                                                                               // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [22:0] id_router_001_src_channel;                                                                                            // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                              // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_001_src2_ready;                                                                                        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	wire          id_router_002_src_endofpacket;                                                                                        // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                              // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                                      // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [106:0] id_router_002_src_data;                                                                                               // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [22:0] id_router_002_src_channel;                                                                                            // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                              // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_demux_001_src3_ready;                                                                                        // timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire          id_router_003_src_endofpacket;                                                                                        // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                              // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                                      // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [106:0] id_router_003_src_data;                                                                                               // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [22:0] id_router_003_src_channel;                                                                                            // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                              // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                                        // timestamp_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_004_src_endofpacket;                                                                                        // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                              // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                                      // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [106:0] id_router_004_src_data;                                                                                               // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [22:0] id_router_004_src_channel;                                                                                            // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                              // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_mux_005_src_endofpacket;                                                                                     // cmd_xbar_mux_005:src_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          cmd_xbar_mux_005_src_valid;                                                                                           // cmd_xbar_mux_005:src_valid -> burst_adapter_001:sink0_valid
	wire          cmd_xbar_mux_005_src_startofpacket;                                                                                   // cmd_xbar_mux_005:src_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [88:0] cmd_xbar_mux_005_src_data;                                                                                            // cmd_xbar_mux_005:src_data -> burst_adapter_001:sink0_data
	wire   [22:0] cmd_xbar_mux_005_src_channel;                                                                                         // cmd_xbar_mux_005:src_channel -> burst_adapter_001:sink0_channel
	wire          cmd_xbar_mux_005_src_ready;                                                                                           // burst_adapter_001:sink0_ready -> cmd_xbar_mux_005:src_ready
	wire          id_router_005_src_endofpacket;                                                                                        // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                              // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                                      // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire   [88:0] id_router_005_src_data;                                                                                               // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [22:0] id_router_005_src_channel;                                                                                            // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                              // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                                        // pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_006_src_endofpacket;                                                                                        // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                              // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                                      // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [106:0] id_router_006_src_data;                                                                                               // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [22:0] id_router_006_src_channel;                                                                                            // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                              // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                                        // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_007_src_endofpacket;                                                                                        // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                              // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                                      // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [106:0] id_router_007_src_data;                                                                                               // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [22:0] id_router_007_src_channel;                                                                                            // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                              // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          width_adapter_003_src_ready;                                                                                          // burst_adapter_002:sink0_ready -> width_adapter_003:out_ready
	wire          id_router_008_src_endofpacket;                                                                                        // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                              // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                                      // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire   [79:0] id_router_008_src_data;                                                                                               // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [22:0] id_router_008_src_channel;                                                                                            // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                              // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_001_src9_ready;                                                                                        // leds_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire          id_router_009_src_endofpacket;                                                                                        // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                              // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                                      // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [106:0] id_router_009_src_data;                                                                                               // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [22:0] id_router_009_src_channel;                                                                                            // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                              // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_001_src10_ready;                                                                                       // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire          id_router_010_src_endofpacket;                                                                                        // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                              // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                                      // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [106:0] id_router_010_src_data;                                                                                               // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [22:0] id_router_010_src_channel;                                                                                            // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                              // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_001_src11_ready;                                                                                       // Switches_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire          id_router_011_src_endofpacket;                                                                                        // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                              // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                                      // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [106:0] id_router_011_src_data;                                                                                               // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [22:0] id_router_011_src_channel;                                                                                            // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                              // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_001_src12_ready;                                                                                       // Keys_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire          id_router_012_src_endofpacket;                                                                                        // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                              // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                                      // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [106:0] id_router_012_src_data;                                                                                               // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [22:0] id_router_012_src_channel;                                                                                            // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                              // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_demux_001_src13_ready;                                                                                       // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	wire          id_router_013_src_endofpacket;                                                                                        // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                              // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                                      // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [106:0] id_router_013_src_data;                                                                                               // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [22:0] id_router_013_src_channel;                                                                                            // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                              // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_001_src14_ready;                                                                                       // audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src14_ready
	wire          id_router_014_src_endofpacket;                                                                                        // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                                              // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                                      // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [106:0] id_router_014_src_data;                                                                                               // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [22:0] id_router_014_src_channel;                                                                                            // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                                              // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_001_src15_ready;                                                                                       // LEDR_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src15_ready
	wire          id_router_015_src_endofpacket;                                                                                        // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                              // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                                      // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [106:0] id_router_015_src_data;                                                                                               // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [22:0] id_router_015_src_channel;                                                                                            // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                              // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_001_src16_ready;                                                                                       // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src16_ready
	wire          id_router_016_src_endofpacket;                                                                                        // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                                              // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                                      // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [106:0] id_router_016_src_data;                                                                                               // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [22:0] id_router_016_src_channel;                                                                                            // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                                              // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          cmd_xbar_demux_001_src17_ready;                                                                                       // hex0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src17_ready
	wire          id_router_017_src_endofpacket;                                                                                        // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                                              // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                                      // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [106:0] id_router_017_src_data;                                                                                               // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [22:0] id_router_017_src_channel;                                                                                            // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                                              // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          cmd_xbar_demux_001_src18_ready;                                                                                       // hex1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src18_ready
	wire          id_router_018_src_endofpacket;                                                                                        // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                                              // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                                      // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [106:0] id_router_018_src_data;                                                                                               // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire   [22:0] id_router_018_src_channel;                                                                                            // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                                              // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          cmd_xbar_demux_001_src19_ready;                                                                                       // hex2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src19_ready
	wire          id_router_019_src_endofpacket;                                                                                        // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire          id_router_019_src_valid;                                                                                              // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire          id_router_019_src_startofpacket;                                                                                      // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [106:0] id_router_019_src_data;                                                                                               // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire   [22:0] id_router_019_src_channel;                                                                                            // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire          id_router_019_src_ready;                                                                                              // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire          cmd_xbar_demux_001_src20_ready;                                                                                       // hex3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src20_ready
	wire          id_router_020_src_endofpacket;                                                                                        // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire          id_router_020_src_valid;                                                                                              // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire          id_router_020_src_startofpacket;                                                                                      // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [106:0] id_router_020_src_data;                                                                                               // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire   [22:0] id_router_020_src_channel;                                                                                            // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire          id_router_020_src_ready;                                                                                              // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire          cmd_xbar_demux_001_src21_ready;                                                                                       // hex4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src21_ready
	wire          id_router_021_src_endofpacket;                                                                                        // id_router_021:src_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire          id_router_021_src_valid;                                                                                              // id_router_021:src_valid -> rsp_xbar_demux_021:sink_valid
	wire          id_router_021_src_startofpacket;                                                                                      // id_router_021:src_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire  [106:0] id_router_021_src_data;                                                                                               // id_router_021:src_data -> rsp_xbar_demux_021:sink_data
	wire   [22:0] id_router_021_src_channel;                                                                                            // id_router_021:src_channel -> rsp_xbar_demux_021:sink_channel
	wire          id_router_021_src_ready;                                                                                              // rsp_xbar_demux_021:sink_ready -> id_router_021:src_ready
	wire          width_adapter_004_src_ready;                                                                                          // burst_adapter_003:sink0_ready -> width_adapter_004:out_ready
	wire          id_router_022_src_endofpacket;                                                                                        // id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire          id_router_022_src_valid;                                                                                              // id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	wire          id_router_022_src_startofpacket;                                                                                      // id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire   [79:0] id_router_022_src_data;                                                                                               // id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	wire   [22:0] id_router_022_src_channel;                                                                                            // id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	wire          id_router_022_src_ready;                                                                                              // rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                                      // cmd_xbar_demux:src1_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                            // cmd_xbar_demux:src1_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                                    // cmd_xbar_demux:src1_startofpacket -> width_adapter:in_startofpacket
	wire  [106:0] cmd_xbar_demux_src1_data;                                                                                             // cmd_xbar_demux:src1_data -> width_adapter:in_data
	wire   [22:0] cmd_xbar_demux_src1_channel;                                                                                          // cmd_xbar_demux:src1_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                            // width_adapter:in_ready -> cmd_xbar_demux:src1_ready
	wire          width_adapter_src_endofpacket;                                                                                        // width_adapter:out_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                              // width_adapter:out_valid -> cmd_xbar_mux_001:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                                      // width_adapter:out_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire   [88:0] width_adapter_src_data;                                                                                               // width_adapter:out_data -> cmd_xbar_mux_001:sink0_data
	wire          width_adapter_src_ready;                                                                                              // cmd_xbar_mux_001:sink0_ready -> width_adapter:out_ready
	wire   [22:0] width_adapter_src_channel;                                                                                            // width_adapter:out_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                                  // cmd_xbar_demux_001:src1_endofpacket -> width_adapter_001:in_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                                        // cmd_xbar_demux_001:src1_valid -> width_adapter_001:in_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                                // cmd_xbar_demux_001:src1_startofpacket -> width_adapter_001:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src1_data;                                                                                         // cmd_xbar_demux_001:src1_data -> width_adapter_001:in_data
	wire   [22:0] cmd_xbar_demux_001_src1_channel;                                                                                      // cmd_xbar_demux_001:src1_channel -> width_adapter_001:in_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                                        // width_adapter_001:in_ready -> cmd_xbar_demux_001:src1_ready
	wire          width_adapter_001_src_endofpacket;                                                                                    // width_adapter_001:out_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          width_adapter_001_src_valid;                                                                                          // width_adapter_001:out_valid -> cmd_xbar_mux_001:sink1_valid
	wire          width_adapter_001_src_startofpacket;                                                                                  // width_adapter_001:out_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire   [88:0] width_adapter_001_src_data;                                                                                           // width_adapter_001:out_data -> cmd_xbar_mux_001:sink1_data
	wire          width_adapter_001_src_ready;                                                                                          // cmd_xbar_mux_001:sink1_ready -> width_adapter_001:out_ready
	wire   [22:0] width_adapter_001_src_channel;                                                                                        // width_adapter_001:out_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                                  // cmd_xbar_demux_001:src5_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                                        // cmd_xbar_demux_001:src5_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                                // cmd_xbar_demux_001:src5_startofpacket -> width_adapter_002:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src5_data;                                                                                         // cmd_xbar_demux_001:src5_data -> width_adapter_002:in_data
	wire   [22:0] cmd_xbar_demux_001_src5_channel;                                                                                      // cmd_xbar_demux_001:src5_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_demux_001_src5_ready;                                                                                        // width_adapter_002:in_ready -> cmd_xbar_demux_001:src5_ready
	wire          width_adapter_002_src_endofpacket;                                                                                    // width_adapter_002:out_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                                          // width_adapter_002:out_valid -> cmd_xbar_mux_005:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                                                  // width_adapter_002:out_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire   [88:0] width_adapter_002_src_data;                                                                                           // width_adapter_002:out_data -> cmd_xbar_mux_005:sink0_data
	wire          width_adapter_002_src_ready;                                                                                          // cmd_xbar_mux_005:sink0_ready -> width_adapter_002:out_ready
	wire   [22:0] width_adapter_002_src_channel;                                                                                        // width_adapter_002:out_channel -> cmd_xbar_mux_005:sink0_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                                                  // cmd_xbar_demux_001:src8_endofpacket -> width_adapter_003:in_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                                        // cmd_xbar_demux_001:src8_valid -> width_adapter_003:in_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                                                // cmd_xbar_demux_001:src8_startofpacket -> width_adapter_003:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src8_data;                                                                                         // cmd_xbar_demux_001:src8_data -> width_adapter_003:in_data
	wire   [22:0] cmd_xbar_demux_001_src8_channel;                                                                                      // cmd_xbar_demux_001:src8_channel -> width_adapter_003:in_channel
	wire          cmd_xbar_demux_001_src8_ready;                                                                                        // width_adapter_003:in_ready -> cmd_xbar_demux_001:src8_ready
	wire          width_adapter_003_src_endofpacket;                                                                                    // width_adapter_003:out_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire          width_adapter_003_src_valid;                                                                                          // width_adapter_003:out_valid -> burst_adapter_002:sink0_valid
	wire          width_adapter_003_src_startofpacket;                                                                                  // width_adapter_003:out_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire   [79:0] width_adapter_003_src_data;                                                                                           // width_adapter_003:out_data -> burst_adapter_002:sink0_data
	wire   [22:0] width_adapter_003_src_channel;                                                                                        // width_adapter_003:out_channel -> burst_adapter_002:sink0_channel
	wire          cmd_xbar_demux_001_src22_endofpacket;                                                                                 // cmd_xbar_demux_001:src22_endofpacket -> width_adapter_004:in_endofpacket
	wire          cmd_xbar_demux_001_src22_valid;                                                                                       // cmd_xbar_demux_001:src22_valid -> width_adapter_004:in_valid
	wire          cmd_xbar_demux_001_src22_startofpacket;                                                                               // cmd_xbar_demux_001:src22_startofpacket -> width_adapter_004:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src22_data;                                                                                        // cmd_xbar_demux_001:src22_data -> width_adapter_004:in_data
	wire   [22:0] cmd_xbar_demux_001_src22_channel;                                                                                     // cmd_xbar_demux_001:src22_channel -> width_adapter_004:in_channel
	wire          cmd_xbar_demux_001_src22_ready;                                                                                       // width_adapter_004:in_ready -> cmd_xbar_demux_001:src22_ready
	wire          width_adapter_004_src_endofpacket;                                                                                    // width_adapter_004:out_endofpacket -> burst_adapter_003:sink0_endofpacket
	wire          width_adapter_004_src_valid;                                                                                          // width_adapter_004:out_valid -> burst_adapter_003:sink0_valid
	wire          width_adapter_004_src_startofpacket;                                                                                  // width_adapter_004:out_startofpacket -> burst_adapter_003:sink0_startofpacket
	wire   [79:0] width_adapter_004_src_data;                                                                                           // width_adapter_004:out_data -> burst_adapter_003:sink0_data
	wire   [22:0] width_adapter_004_src_channel;                                                                                        // width_adapter_004:out_channel -> burst_adapter_003:sink0_channel
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                                  // rsp_xbar_demux_001:src0_endofpacket -> width_adapter_005:in_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                                        // rsp_xbar_demux_001:src0_valid -> width_adapter_005:in_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                                // rsp_xbar_demux_001:src0_startofpacket -> width_adapter_005:in_startofpacket
	wire   [88:0] rsp_xbar_demux_001_src0_data;                                                                                         // rsp_xbar_demux_001:src0_data -> width_adapter_005:in_data
	wire   [22:0] rsp_xbar_demux_001_src0_channel;                                                                                      // rsp_xbar_demux_001:src0_channel -> width_adapter_005:in_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                                        // width_adapter_005:in_ready -> rsp_xbar_demux_001:src0_ready
	wire          width_adapter_005_src_endofpacket;                                                                                    // width_adapter_005:out_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          width_adapter_005_src_valid;                                                                                          // width_adapter_005:out_valid -> rsp_xbar_mux:sink1_valid
	wire          width_adapter_005_src_startofpacket;                                                                                  // width_adapter_005:out_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [106:0] width_adapter_005_src_data;                                                                                           // width_adapter_005:out_data -> rsp_xbar_mux:sink1_data
	wire          width_adapter_005_src_ready;                                                                                          // rsp_xbar_mux:sink1_ready -> width_adapter_005:out_ready
	wire   [22:0] width_adapter_005_src_channel;                                                                                        // width_adapter_005:out_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                                  // rsp_xbar_demux_001:src1_endofpacket -> width_adapter_006:in_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                                        // rsp_xbar_demux_001:src1_valid -> width_adapter_006:in_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                                // rsp_xbar_demux_001:src1_startofpacket -> width_adapter_006:in_startofpacket
	wire   [88:0] rsp_xbar_demux_001_src1_data;                                                                                         // rsp_xbar_demux_001:src1_data -> width_adapter_006:in_data
	wire   [22:0] rsp_xbar_demux_001_src1_channel;                                                                                      // rsp_xbar_demux_001:src1_channel -> width_adapter_006:in_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                                        // width_adapter_006:in_ready -> rsp_xbar_demux_001:src1_ready
	wire          width_adapter_006_src_endofpacket;                                                                                    // width_adapter_006:out_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          width_adapter_006_src_valid;                                                                                          // width_adapter_006:out_valid -> rsp_xbar_mux_001:sink1_valid
	wire          width_adapter_006_src_startofpacket;                                                                                  // width_adapter_006:out_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [106:0] width_adapter_006_src_data;                                                                                           // width_adapter_006:out_data -> rsp_xbar_mux_001:sink1_data
	wire          width_adapter_006_src_ready;                                                                                          // rsp_xbar_mux_001:sink1_ready -> width_adapter_006:out_ready
	wire   [22:0] width_adapter_006_src_channel;                                                                                        // width_adapter_006:out_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                                  // rsp_xbar_demux_005:src0_endofpacket -> width_adapter_007:in_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                                        // rsp_xbar_demux_005:src0_valid -> width_adapter_007:in_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                                // rsp_xbar_demux_005:src0_startofpacket -> width_adapter_007:in_startofpacket
	wire   [88:0] rsp_xbar_demux_005_src0_data;                                                                                         // rsp_xbar_demux_005:src0_data -> width_adapter_007:in_data
	wire   [22:0] rsp_xbar_demux_005_src0_channel;                                                                                      // rsp_xbar_demux_005:src0_channel -> width_adapter_007:in_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                                        // width_adapter_007:in_ready -> rsp_xbar_demux_005:src0_ready
	wire          width_adapter_007_src_endofpacket;                                                                                    // width_adapter_007:out_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          width_adapter_007_src_valid;                                                                                          // width_adapter_007:out_valid -> rsp_xbar_mux_001:sink5_valid
	wire          width_adapter_007_src_startofpacket;                                                                                  // width_adapter_007:out_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [106:0] width_adapter_007_src_data;                                                                                           // width_adapter_007:out_data -> rsp_xbar_mux_001:sink5_data
	wire          width_adapter_007_src_ready;                                                                                          // rsp_xbar_mux_001:sink5_ready -> width_adapter_007:out_ready
	wire   [22:0] width_adapter_007_src_channel;                                                                                        // width_adapter_007:out_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                                  // rsp_xbar_demux_008:src0_endofpacket -> width_adapter_008:in_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                                        // rsp_xbar_demux_008:src0_valid -> width_adapter_008:in_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                                // rsp_xbar_demux_008:src0_startofpacket -> width_adapter_008:in_startofpacket
	wire   [79:0] rsp_xbar_demux_008_src0_data;                                                                                         // rsp_xbar_demux_008:src0_data -> width_adapter_008:in_data
	wire   [22:0] rsp_xbar_demux_008_src0_channel;                                                                                      // rsp_xbar_demux_008:src0_channel -> width_adapter_008:in_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                                        // width_adapter_008:in_ready -> rsp_xbar_demux_008:src0_ready
	wire          width_adapter_008_src_endofpacket;                                                                                    // width_adapter_008:out_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          width_adapter_008_src_valid;                                                                                          // width_adapter_008:out_valid -> rsp_xbar_mux_001:sink8_valid
	wire          width_adapter_008_src_startofpacket;                                                                                  // width_adapter_008:out_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [106:0] width_adapter_008_src_data;                                                                                           // width_adapter_008:out_data -> rsp_xbar_mux_001:sink8_data
	wire          width_adapter_008_src_ready;                                                                                          // rsp_xbar_mux_001:sink8_ready -> width_adapter_008:out_ready
	wire   [22:0] width_adapter_008_src_channel;                                                                                        // width_adapter_008:out_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_022_src0_endofpacket;                                                                                  // rsp_xbar_demux_022:src0_endofpacket -> width_adapter_009:in_endofpacket
	wire          rsp_xbar_demux_022_src0_valid;                                                                                        // rsp_xbar_demux_022:src0_valid -> width_adapter_009:in_valid
	wire          rsp_xbar_demux_022_src0_startofpacket;                                                                                // rsp_xbar_demux_022:src0_startofpacket -> width_adapter_009:in_startofpacket
	wire   [79:0] rsp_xbar_demux_022_src0_data;                                                                                         // rsp_xbar_demux_022:src0_data -> width_adapter_009:in_data
	wire   [22:0] rsp_xbar_demux_022_src0_channel;                                                                                      // rsp_xbar_demux_022:src0_channel -> width_adapter_009:in_channel
	wire          rsp_xbar_demux_022_src0_ready;                                                                                        // width_adapter_009:in_ready -> rsp_xbar_demux_022:src0_ready
	wire          width_adapter_009_src_endofpacket;                                                                                    // width_adapter_009:out_endofpacket -> rsp_xbar_mux_001:sink22_endofpacket
	wire          width_adapter_009_src_valid;                                                                                          // width_adapter_009:out_valid -> rsp_xbar_mux_001:sink22_valid
	wire          width_adapter_009_src_startofpacket;                                                                                  // width_adapter_009:out_startofpacket -> rsp_xbar_mux_001:sink22_startofpacket
	wire  [106:0] width_adapter_009_src_data;                                                                                           // width_adapter_009:out_data -> rsp_xbar_mux_001:sink22_data
	wire          width_adapter_009_src_ready;                                                                                          // rsp_xbar_mux_001:sink22_ready -> width_adapter_009:out_ready
	wire   [22:0] width_adapter_009_src_channel;                                                                                        // width_adapter_009:out_channel -> rsp_xbar_mux_001:sink22_channel
	wire   [22:0] limiter_cmd_valid_data;                                                                                               // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [22:0] limiter_001_cmd_valid_data;                                                                                           // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                                             // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                                             // timer:irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                                             // timestamp:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                                                             // audio:irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                                                             // Keys:irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                                                                             // Switches:irq -> irq_mapper:receiver5_irq
	wire          irq_mapper_receiver6_irq;                                                                                             // ps2_0:irq -> irq_mapper:receiver6_irq
	wire   [31:0] nios2_processor_d_irq_irq;                                                                                            // irq_mapper:sender_irq -> nios2_processor:d_irq

	nios_system_nios2_processor nios2_processor (
		.clk                                   (clocks_sys_clk_clk),                                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                                //                   reset_n.reset_n
		.d_address                             (nios2_processor_data_master_address),                                            //               data_master.address
		.d_byteenable                          (nios2_processor_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (nios2_processor_data_master_read),                                               //                          .read
		.d_readdata                            (nios2_processor_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (nios2_processor_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (nios2_processor_data_master_write),                                              //                          .write
		.d_writedata                           (nios2_processor_data_master_writedata),                                          //                          .writedata
		.d_readdatavalid                       (nios2_processor_data_master_readdatavalid),                                      //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_processor_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (nios2_processor_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (nios2_processor_instruction_master_read),                                        //                          .read
		.i_readdata                            (nios2_processor_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (nios2_processor_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (nios2_processor_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (nios2_processor_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_processor_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                                // custom_instruction_master.readra
	);

	nios_system_jtag_uart jtag_uart (
		.clk            (clocks_sys_clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                //               irq.irq
	);

	nios_system_sdram sdram (
		.clk            (clocks_sys_clk_clk),                                    //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                       // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_wire_dq),                                         //      .export
		.zs_dqm         (sdram_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_wire_we_n)                                        //      .export
	);

	nios_system_timer timer (
		.clk        (clocks_sys_clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    // reset.reset_n
		.address    (timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                            //   irq.irq
	);

	nios_system_clocks clocks (
		.CLOCK_50    (clk_clk),                            //       clk_in_primary.clk
		.reset       (rst_controller_001_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (clocks_sys_clk_clk),                 //              sys_clk.clk
		.sys_reset_n (),                                   //        sys_clk_reset.reset_n
		.SDRAM_CLK   (sdram_clk_clk),                      //            sdram_clk.clk
		.VGA_CLK     (clocks_vga_clk_clk)                  //              vga_clk.clk
	);

	nios_system_timer timestamp (
		.clk        (clocks_sys_clk_clk),                                     //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        // reset.reset_n
		.address    (timestamp_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timestamp_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timestamp_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timestamp_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timestamp_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                                //   irq.irq
	);

	nios_system_pixel_buffer pixel_buffer (
		.clk           (clocks_sys_clk_clk),                                                          //        clock_reset.clk
		.reset         (rst_controller_reset_out_reset),                                              //  clock_reset_reset.reset
		.SRAM_DQ       (sram_interface_DQ),                                                           // external_interface.export
		.SRAM_ADDR     (sram_interface_ADDR),                                                         //                   .export
		.SRAM_LB_N     (sram_interface_LB_N),                                                         //                   .export
		.SRAM_UB_N     (sram_interface_UB_N),                                                         //                   .export
		.SRAM_CE_N     (sram_interface_CE_N),                                                         //                   .export
		.SRAM_OE_N     (sram_interface_OE_N),                                                         //                   .export
		.SRAM_WE_N     (sram_interface_WE_N),                                                         //                   .export
		.address       (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address),       //  avalon_sram_slave.address
		.byteenable    (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.read          (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read),          //                   .read
		.write         (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write),         //                   .write
		.writedata     (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.readdata      (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.readdatavalid (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid)  //                   .readdatavalid
	);

	nios_system_pixel_buffer_dma_0 pixel_buffer_dma_0 (
		.clk                  (clocks_sys_clk_clk),                                                                //             clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                                                    //       clock_reset_reset.reset
		.master_readdatavalid (pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid),                          // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest),                            //                        .waitrequest
		.master_address       (pixel_buffer_dma_0_avalon_pixel_dma_master_address),                                //                        .address
		.master_arbiterlock   (pixel_buffer_dma_0_avalon_pixel_dma_master_lock),                                   //                        .lock
		.master_read          (pixel_buffer_dma_0_avalon_pixel_dma_master_read),                                   //                        .read
		.master_readdata      (pixel_buffer_dma_0_avalon_pixel_dma_master_readdata),                               //                        .readdata
		.slave_address        (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_address),    //    avalon_control_slave.address
		.slave_byteenable     (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_byteenable), //                        .byteenable
		.slave_read           (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_read),       //                        .read
		.slave_write          (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_write),      //                        .write
		.slave_writedata      (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_writedata),  //                        .writedata
		.slave_readdata       (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_readdata),   //                        .readdata
		.stream_ready         (pixel_buffer_dma_0_avalon_pixel_source_ready),                                      //     avalon_pixel_source.ready
		.stream_startofpacket (pixel_buffer_dma_0_avalon_pixel_source_startofpacket),                              //                        .startofpacket
		.stream_endofpacket   (pixel_buffer_dma_0_avalon_pixel_source_endofpacket),                                //                        .endofpacket
		.stream_valid         (pixel_buffer_dma_0_avalon_pixel_source_valid),                                      //                        .valid
		.stream_data          (pixel_buffer_dma_0_avalon_pixel_source_data)                                        //                        .data
	);

	nios_system_rgb_resampler rgb_resampler (
		.clk                      (clocks_sys_clk_clk),                                   //       clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                       // clock_reset_reset.reset
		.stream_in_startofpacket  (pixel_buffer_dma_0_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (pixel_buffer_dma_0_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (pixel_buffer_dma_0_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (pixel_buffer_dma_0_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (pixel_buffer_dma_0_avalon_pixel_source_data),          //                  .data
		.stream_out_ready         (rgb_resampler_avalon_rgb_source_ready),                // avalon_rgb_source.ready
		.stream_out_startofpacket (rgb_resampler_avalon_rgb_source_startofpacket),        //                  .startofpacket
		.stream_out_endofpacket   (rgb_resampler_avalon_rgb_source_endofpacket),          //                  .endofpacket
		.stream_out_valid         (rgb_resampler_avalon_rgb_source_valid),                //                  .valid
		.stream_out_data          (rgb_resampler_avalon_rgb_source_data)                  //                  .data
	);

	nios_system_scaler scaler (
		.clk                      (clocks_sys_clk_clk),                            //          clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                //    clock_reset_reset.reset
		.stream_in_startofpacket  (rgb_resampler_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (rgb_resampler_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (rgb_resampler_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (rgb_resampler_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (rgb_resampler_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (scaler_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (scaler_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (scaler_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (scaler_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (scaler_avalon_scaler_source_data)               //                     .data
	);

	nios_system_video_fifo video_fifo (
		.clk_stream_in            (clocks_sys_clk_clk),                                //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                    //   clock_stream_in_reset.reset
		.clk_stream_out           (clocks_vga_clk_clk),                                //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),                //  clock_stream_out_reset.reset
		.stream_in_ready          (alpha_blender_avalon_blended_source_ready),         //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (alpha_blender_avalon_blended_source_startofpacket), //                        .startofpacket
		.stream_in_endofpacket    (alpha_blender_avalon_blended_source_endofpacket),   //                        .endofpacket
		.stream_in_valid          (alpha_blender_avalon_blended_source_valid),         //                        .valid
		.stream_in_data           (alpha_blender_avalon_blended_source_data),          //                        .data
		.stream_out_ready         (video_fifo_avalon_dc_buffer_source_ready),          // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (video_fifo_avalon_dc_buffer_source_startofpacket),  //                        .startofpacket
		.stream_out_endofpacket   (video_fifo_avalon_dc_buffer_source_endofpacket),    //                        .endofpacket
		.stream_out_valid         (video_fifo_avalon_dc_buffer_source_valid),          //                        .valid
		.stream_out_data          (video_fifo_avalon_dc_buffer_source_data)            //                        .data
	);

	nios_system_vga_controller vga_controller (
		.clk           (clocks_vga_clk_clk),                               //        clock_reset.clk
		.reset         (rst_controller_002_reset_out_reset),               //  clock_reset_reset.reset
		.data          (video_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (video_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (video_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_extern_CLK),                                   // external_interface.export
		.VGA_HS        (vga_extern_HS),                                    //                   .export
		.VGA_VS        (vga_extern_VS),                                    //                   .export
		.VGA_BLANK     (vga_extern_BLANK),                                 //                   .export
		.VGA_SYNC      (vga_extern_SYNC),                                  //                   .export
		.VGA_R         (vga_extern_R),                                     //                   .export
		.VGA_G         (vga_extern_G),                                     //                   .export
		.VGA_B         (vga_extern_B)                                      //                   .export
	);

	nios_system_char_drawer char_drawer (
		.clk                  (clocks_sys_clk_clk),                                                              //               clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                                                  //         clock_reset_reset.reset
		.ctrl_address         (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable), //                          .byteenable
		.ctrl_chipselect      (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect), //                          .chipselect
		.ctrl_read            (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_read),       //                          .read
		.ctrl_write           (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_write),      //                          .write
		.ctrl_writedata       (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata),  //                          .writedata
		.ctrl_readdata        (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata),   //                          .readdata
		.buf_byteenable       (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect),  //                          .chipselect
		.buf_read             (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read),        //                          .read
		.buf_write            (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write),       //                          .write
		.buf_writedata        (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.buf_readdata         (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.buf_waitrequest      (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.buf_address          (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address),     //                          .address
		.stream_ready         (char_drawer_avalon_char_source_ready),                                            //        avalon_char_source.ready
		.stream_startofpacket (char_drawer_avalon_char_source_startofpacket),                                    //                          .startofpacket
		.stream_endofpacket   (char_drawer_avalon_char_source_endofpacket),                                      //                          .endofpacket
		.stream_valid         (char_drawer_avalon_char_source_valid),                                            //                          .valid
		.stream_data          (char_drawer_avalon_char_source_data)                                              //                          .data
	);

	nios_system_alpha_blender alpha_blender (
		.clk                      (clocks_sys_clk_clk),                                //            clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                    //      clock_reset_reset.reset
		.foreground_data          (char_drawer_avalon_char_source_data),               // avalon_foreground_sink.data
		.foreground_startofpacket (char_drawer_avalon_char_source_startofpacket),      //                       .startofpacket
		.foreground_endofpacket   (char_drawer_avalon_char_source_endofpacket),        //                       .endofpacket
		.foreground_valid         (char_drawer_avalon_char_source_valid),              //                       .valid
		.foreground_ready         (char_drawer_avalon_char_source_ready),              //                       .ready
		.background_data          (scaler_avalon_scaler_source_data),                  // avalon_background_sink.data
		.background_startofpacket (scaler_avalon_scaler_source_startofpacket),         //                       .startofpacket
		.background_endofpacket   (scaler_avalon_scaler_source_endofpacket),           //                       .endofpacket
		.background_valid         (scaler_avalon_scaler_source_valid),                 //                       .valid
		.background_ready         (scaler_avalon_scaler_source_ready),                 //                       .ready
		.output_ready             (alpha_blender_avalon_blended_source_ready),         //  avalon_blended_source.ready
		.output_data              (alpha_blender_avalon_blended_source_data),          //                       .data
		.output_startofpacket     (alpha_blender_avalon_blended_source_startofpacket), //                       .startofpacket
		.output_endofpacket       (alpha_blender_avalon_blended_source_endofpacket),   //                       .endofpacket
		.output_valid             (alpha_blender_avalon_blended_source_valid)          //                       .valid
	);

	nios_system_leds leds (
		.clk        (clocks_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (leds_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~leds_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (leds_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (leds_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (leds_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (leds_export)                                        // external_connection.export
	);

	Altera_UP_SD_Card_Avalon_Interface sd_card (
		.i_avalon_chip_select (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_address),     //                    .address
		.i_avalon_read        (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_read),        //                    .read
		.i_avalon_write       (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_write),       //                    .write
		.i_avalon_byteenable  (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable),  //                    .byteenable
		.i_avalon_writedata   (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata),   //                    .writedata
		.o_avalon_readdata    (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata),    //                    .readdata
		.o_avalon_waitrequest (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest), //                    .waitrequest
		.i_clock              (clocks_sys_clk_clk),                                                     //          clock_sink.clk
		.i_reset_n            (~rst_controller_reset_out_reset),                                        //    clock_sink_reset.reset_n
		.b_SD_cmd             (sd_card_b_SD_cmd),                                                       //         conduit_end.export
		.b_SD_dat             (sd_card_b_SD_dat),                                                       //                    .export
		.b_SD_dat3            (sd_card_b_SD_dat3),                                                      //                    .export
		.o_SD_clock           (sd_card_o_SD_clock)                                                      //                    .export
	);

	nios_system_Keys keys (
		.clk        (clocks_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (keys_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~keys_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (keys_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (keys_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (keys_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (keys_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                           //                 irq.irq
	);

	nios_system_Switches switches (
		.clk        (clocks_sys_clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (switches_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~switches_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (switches_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (switches_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (switches_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (switches_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                               //                 irq.irq
	);

	nios_system_audio_and_video_config_0 audio_and_video_config_0 (
		.clk         (clocks_sys_clk_clk),                                                                         //            clock_reset.clk
		.reset       (rst_controller_003_reset_out_reset),                                                         //      clock_reset_reset.reset
		.address     (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_address),     // avalon_av_config_slave.address
		.byteenable  (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),  //                       .byteenable
		.read        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_read),        //                       .read
		.write       (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_write),       //                       .write
		.writedata   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),   //                       .writedata
		.readdata    (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),    //                       .readdata
		.waitrequest (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest), //                       .waitrequest
		.I2C_SDAT    (audio_and_video_config_SDAT),                                                                //     external_interface.export
		.I2C_SCLK    (audio_and_video_config_SCLK)                                                                 //                       .export
	);

	nios_system_up_clocks_0 up_clocks_0 (
		.CLOCK_50    (clocks_sys_clk_clk),                 //       clk_in_primary.clk
		.reset       (rst_controller_003_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (),                                   //              sys_clk.clk
		.sys_reset_n (),                                   //        sys_clk_reset.reset_n
		.CLOCK_27    (clk_in_secondary_clk),               //     clk_in_secondary.clk
		.AUD_CLK     (audio_clk_clk)                       //            audio_clk.clk
	);

	nios_system_audio audio (
		.clk         (clocks_sys_clk_clk),                                                 //        clock_reset.clk
		.reset       (rst_controller_003_reset_out_reset),                                 //  clock_reset_reset.reset
		.address     (audio_avalon_audio_slave_translator_avalon_anti_slave_0_address),    // avalon_audio_slave.address
		.chipselect  (audio_avalon_audio_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.read        (audio_avalon_audio_slave_translator_avalon_anti_slave_0_read),       //                   .read
		.write       (audio_avalon_audio_slave_translator_avalon_anti_slave_0_write),      //                   .write
		.writedata   (audio_avalon_audio_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.readdata    (audio_avalon_audio_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.irq         (irq_mapper_receiver3_irq),                                           //          interrupt.irq
		.AUD_ADCDAT  (audio_ADCDAT),                                                       // external_interface.export
		.AUD_ADCLRCK (audio_ADCLRCK),                                                      //                   .export
		.AUD_BCLK    (audio_BCLK),                                                         //                   .export
		.AUD_DACDAT  (audio_DACDAT),                                                       //                   .export
		.AUD_DACLRCK (audio_DACLRCK)                                                       //                   .export
	);

	nios_system_LEDR ledr (
		.clk        (clocks_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (ledr_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ledr_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ledr_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ledr_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ledr_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ledrs_export)                                       // external_connection.export
	);

	nios_system_ps2_0 ps2_0 (
		.clk         (clocks_sys_clk_clk),                                                //        clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                    //  clock_reset_reset.reset
		.address     (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_address),     //   avalon_ps2_slave.address
		.chipselect  (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_chipselect),  //                   .chipselect
		.byteenable  (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_byteenable),  //                   .byteenable
		.read        (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_read),        //                   .read
		.write       (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_write),       //                   .write
		.writedata   (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.readdata    (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.waitrequest (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.irq         (irq_mapper_receiver6_irq),                                          //          interrupt.irq
		.PS2_CLK     (ps2_0_external_interface_CLK),                                      // external_interface.export
		.PS2_DAT     (ps2_0_external_interface_DAT)                                       //                   .export
	);

	nios_system_leds hex0 (
		.clk        (clocks_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (hex0_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex0_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex0_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex0_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex0_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex0_ex_export)                                     // external_connection.export
	);

	nios_system_leds hex1 (
		.clk        (clocks_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (hex1_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex1_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex1_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex1_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex1_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex1_ex_export)                                     // external_connection.export
	);

	nios_system_leds hex2 (
		.clk        (clocks_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (hex2_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex2_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex2_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex2_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex2_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex2_ex_export)                                     // external_connection.export
	);

	nios_system_leds hex3 (
		.clk        (clocks_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (hex3_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex3_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex3_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex3_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex3_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex3_ex_export)                                     // external_connection.export
	);

	nios_system_leds hex4 (
		.clk        (clocks_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (hex4_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex4_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex4_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex4_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex4_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex4_ex_export)                                     // external_connection.export
	);

	nios_system_character_lcd_0 character_lcd_0 (
		.clk         (clocks_sys_clk_clk),                                                          //        clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                              //  clock_reset_reset.reset
		.address     (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address),     //   avalon_lcd_slave.address
		.chipselect  (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),  //                   .chipselect
		.read        (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read),        //                   .read
		.write       (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write),       //                   .write
		.writedata   (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.readdata    (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.waitrequest (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.LCD_DATA    (character_lcd_0_external_interface_DATA),                                     // external_interface.export
		.LCD_ON      (character_lcd_0_external_interface_ON),                                       //                   .export
		.LCD_BLON    (character_lcd_0_external_interface_BLON),                                     //                   .export
		.LCD_EN      (character_lcd_0_external_interface_EN),                                       //                   .export
		.LCD_RS      (character_lcd_0_external_interface_RS),                                       //                   .export
		.LCD_RW      (character_lcd_0_external_interface_RW)                                        //                   .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_processor_instruction_master_translator (
		.clk                   (clocks_sys_clk_clk),                                                                    //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                        //                     reset.reset
		.uav_address           (nios2_processor_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_processor_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_processor_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_processor_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_processor_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_processor_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_processor_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_processor_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_processor_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_processor_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_processor_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_processor_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_processor_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (nios2_processor_instruction_master_read),                                               //                          .read
		.av_readdata           (nios2_processor_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_processor_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                                  //               (terminated)
		.av_byteenable         (4'b1111),                                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                  //               (terminated)
		.av_begintransfer      (1'b0),                                                                                  //               (terminated)
		.av_chipselect         (1'b0),                                                                                  //               (terminated)
		.av_write              (1'b0),                                                                                  //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                                  //               (terminated)
		.av_lock               (1'b0),                                                                                  //               (terminated)
		.av_debugaccess        (1'b0),                                                                                  //               (terminated)
		.uav_clken             (),                                                                                      //               (terminated)
		.av_clken              (1'b1)                                                                                   //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_processor_data_master_translator (
		.clk                   (clocks_sys_clk_clk),                                                             //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                     reset.reset
		.uav_address           (nios2_processor_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_processor_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_processor_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_processor_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_processor_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_processor_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_processor_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_processor_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_processor_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_processor_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_processor_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_processor_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_processor_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (nios2_processor_data_master_byteenable),                                         //                          .byteenable
		.av_read               (nios2_processor_data_master_read),                                               //                          .read
		.av_readdata           (nios2_processor_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_processor_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (nios2_processor_data_master_write),                                              //                          .write
		.av_writedata          (nios2_processor_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (nios2_processor_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                           //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                           //               (terminated)
		.av_begintransfer      (1'b0),                                                                           //               (terminated)
		.av_chipselect         (1'b0),                                                                           //               (terminated)
		.av_lock               (1'b0),                                                                           //               (terminated)
		.uav_clken             (),                                                                               //               (terminated)
		.av_clken              (1'b1)                                                                            //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) pixel_buffer_dma_0_avalon_pixel_dma_master_translator (
		.clk                   (clocks_sys_clk_clk),                                                                            //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                //                     reset.reset
		.uav_address           (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (pixel_buffer_dma_0_avalon_pixel_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest),                                        //                          .waitrequest
		.av_read               (pixel_buffer_dma_0_avalon_pixel_dma_master_read),                                               //                          .read
		.av_readdata           (pixel_buffer_dma_0_avalon_pixel_dma_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid),                                      //                          .readdatavalid
		.av_lock               (pixel_buffer_dma_0_avalon_pixel_dma_master_lock),                                               //                          .lock
		.av_burstcount         (1'b1),                                                                                          //               (terminated)
		.av_byteenable         (2'b11),                                                                                         //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                          //               (terminated)
		.av_begintransfer      (1'b0),                                                                                          //               (terminated)
		.av_chipselect         (1'b0),                                                                                          //               (terminated)
		.av_write              (1'b0),                                                                                          //               (terminated)
		.av_writedata          (16'b0000000000000000),                                                                          //               (terminated)
		.av_debugaccess        (1'b0),                                                                                          //               (terminated)
		.uav_clken             (),                                                                                              //               (terminated)
		.av_clken              (1'b1)                                                                                           //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_processor_jtag_debug_module_translator (
		.clk                   (clocks_sys_clk_clk),                                                                           //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                               //                    reset.reset
		.uav_address           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                                             //              (terminated)
		.av_burstcount         (),                                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                                             //              (terminated)
		.av_lock               (),                                                                                             //              (terminated)
		.av_clken              (),                                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_byteenable         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address           (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                    //              (terminated)
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_byteenable         (),                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timestamp_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timestamp_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timestamp_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timestamp_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timestamp_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timestamp_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pixel_buffer_avalon_sram_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer      (),                                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                                          //              (terminated)
		.av_burstcount         (),                                                                                          //              (terminated)
		.av_waitrequest        (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                                          //              (terminated)
		.av_lock               (),                                                                                          //              (terminated)
		.av_chipselect         (),                                                                                          //              (terminated)
		.av_clken              (),                                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                                      //              (terminated)
		.av_debugaccess        (),                                                                                          //              (terminated)
		.av_outputenable       ()                                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pixel_buffer_dma_0_avalon_control_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                     //                    reset.reset
		.uav_address           (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer      (),                                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                                   //              (terminated)
		.av_lock               (),                                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                                   //              (terminated)
		.av_clken              (),                                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) char_drawer_avalon_char_control_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                   //                    reset.reset
		.uav_address           (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                                 //              (terminated)
		.av_lock               (),                                                                                                 //              (terminated)
		.av_clken              (),                                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) char_drawer_avalon_char_buffer_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                  //                    reset.reset
		.uav_address           (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                                //              (terminated)
		.av_burstcount         (),                                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                                //              (terminated)
		.av_lock               (),                                                                                                //              (terminated)
		.av_clken              (),                                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                                //              (terminated)
		.av_outputenable       ()                                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) leds_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (leds_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (leds_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (leds_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (leds_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (leds_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (leds_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (leds_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (leds_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_card_avalon_sdcard_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switches_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address           (switches_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (switches_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (switches_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (switches_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (switches_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (switches_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (switches_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (switches_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (switches_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (switches_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (switches_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (switches_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (switches_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (switches_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_byteenable         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) keys_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (keys_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (keys_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (keys_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (keys_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (keys_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (keys_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (keys_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (keys_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (keys_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (keys_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (keys_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (keys_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (keys_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (keys_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (keys_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (keys_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_and_video_config_0_avalon_av_config_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                                         //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                                         //                    reset.reset
		.uav_address           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                                                           //              (terminated)
		.av_burstcount         (),                                                                                                           //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                                       //              (terminated)
		.av_writebyteenable    (),                                                                                                           //              (terminated)
		.av_lock               (),                                                                                                           //              (terminated)
		.av_chipselect         (),                                                                                                           //              (terminated)
		.av_clken              (),                                                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                                                       //              (terminated)
		.av_debugaccess        (),                                                                                                           //              (terminated)
		.av_outputenable       ()                                                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_avalon_audio_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                  //                    reset.reset
		.uav_address           (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (audio_avalon_audio_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (audio_avalon_audio_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (audio_avalon_audio_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (audio_avalon_audio_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (audio_avalon_audio_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (audio_avalon_audio_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                                    //              (terminated)
		.av_burstcount         (),                                                                                    //              (terminated)
		.av_byteenable         (),                                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                    //              (terminated)
		.av_lock               (),                                                                                    //              (terminated)
		.av_clken              (),                                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                                //              (terminated)
		.av_debugaccess        (),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ledr_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ledr_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ledr_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ledr_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ledr_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (ledr_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ps2_0_avalon_ps2_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address           (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex0_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (hex0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (hex0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (hex0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (hex0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (hex0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (hex0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (hex0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (hex0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (hex0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (hex0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (hex0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (hex0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (hex0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (hex0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex1_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (hex1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (hex1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (hex1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (hex1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (hex1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (hex1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (hex1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (hex1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (hex1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (hex1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (hex1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (hex1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (hex1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (hex1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex2_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (hex2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (hex2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (hex2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (hex2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (hex2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (hex2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (hex2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (hex2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (hex2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (hex2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (hex2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (hex2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (hex2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (hex2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex3_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (hex3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (hex3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (hex3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (hex3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (hex3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (hex3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (hex3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (hex3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (hex3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (hex3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (hex3_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (hex3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (hex3_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (hex3_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex4_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (hex4_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (hex4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (hex4_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (hex4_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (hex4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (hex4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (hex4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (hex4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (hex4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (hex4_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (hex4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (hex4_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (hex4_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (hex4_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (hex4_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (hex4_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) character_lcd_0_avalon_lcd_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                              //                    reset.reset
		.uav_address           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                                            //              (terminated)
		.av_burstcount         (),                                                                                            //              (terminated)
		.av_byteenable         (),                                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                                            //              (terminated)
		.av_lock               (),                                                                                            //              (terminated)
		.av_clken              (),                                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                                        //              (terminated)
		.av_debugaccess        (),                                                                                            //              (terminated)
		.av_outputenable       ()                                                                                             //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (86),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (23),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) nios2_processor_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clocks_sys_clk_clk),                                                                             //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.av_address       (nios2_processor_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_processor_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_processor_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_processor_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_processor_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_processor_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_processor_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_processor_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_processor_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_processor_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_processor_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                                          //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                                           //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                                        //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                                  //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                                    //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                                           //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (86),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (23),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) nios2_processor_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clocks_sys_clk_clk),                                                                      //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.av_address       (nios2_processor_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_processor_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_processor_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_processor_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_processor_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_processor_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_processor_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_processor_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_processor_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_processor_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_processor_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                               //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                                //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                             //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                       //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                         //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                                //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_BEGIN_BURST           (68),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (73),
		.PKT_SRC_ID_L              (69),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (74),
		.PKT_THREAD_ID_H           (79),
		.PKT_THREAD_ID_L           (79),
		.PKT_CACHE_H               (86),
		.PKT_CACHE_L               (83),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (23),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent (
		.clk              (clocks_sys_clk_clk),                                                                                     //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                                         // clk_reset.reset
		.av_address       (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_005_src1_valid),                                                                          //        rp.valid
		.rp_data          (rsp_xbar_demux_005_src1_data),                                                                           //          .data
		.rp_channel       (rsp_xbar_demux_005_src1_channel),                                                                        //          .channel
		.rp_startofpacket (rsp_xbar_demux_005_src1_startofpacket),                                                                  //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_005_src1_endofpacket),                                                                    //          .endofpacket
		.rp_ready         (rsp_xbar_demux_005_src1_ready)                                                                           //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                         //       clk_reset.reset
		.m0_address              (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                                 //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                               //                .channel
		.rf_sink_ready           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                         // clk_reset.reset
		.in_data           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (68),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (73),
		.PKT_SRC_ID_L              (69),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (74),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                   //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                   //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                    //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                             //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                 //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src2_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src2_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src2_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src2_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src2_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src2_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                               //                .channel
		.rf_sink_ready           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timestamp_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                   //                .channel
		.rf_sink_ready           (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (68),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (73),
		.PKT_SRC_ID_L              (69),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (74),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                                     //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                                     //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                                      //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                               //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                                   //                .channel
		.rf_sink_ready           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                               //       clk_reset.reset
		.m0_address              (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                                              //                .channel
		.rf_sink_ready           (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                               // clk_reset.reset
		.in_data           (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                                         // (terminated)
		.csr_readdata      (),                                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                         // (terminated)
		.almost_full_data  (),                                                                                                             // (terminated)
		.almost_empty_data (),                                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                                         // (terminated)
		.out_empty         (),                                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                                         // (terminated)
		.out_error         (),                                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                                         // (terminated)
		.out_channel       ()                                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                             //       clk_reset.reset
		.m0_address              (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                                            //                .channel
		.rf_sink_ready           (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                             // clk_reset.reset
		.in_data           (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                                       // (terminated)
		.csr_readdata      (),                                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                       // (terminated)
		.almost_full_data  (),                                                                                                           // (terminated)
		.almost_empty_data (),                                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                                       // (terminated)
		.out_empty         (),                                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                                       // (terminated)
		.out_error         (),                                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                                       // (terminated)
		.out_channel       ()                                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (59),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (64),
		.PKT_SRC_ID_L              (60),
		.PKT_DEST_ID_H             (69),
		.PKT_DEST_ID_L             (65),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (73),
		.PKT_PROTECTION_L          (71),
		.PKT_RESPONSE_STATUS_H     (79),
		.PKT_RESPONSE_STATUS_L     (78),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (80),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                            //       clk_reset.reset
		.m0_address              (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                                           //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                                           //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                                            //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                                                   //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                                                     //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                                         //                .channel
		.rf_sink_ready           (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (81),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                            // clk_reset.reset
		.in_data           (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                                      // (terminated)
		.csr_readdata      (),                                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                      // (terminated)
		.almost_full_data  (),                                                                                                          // (terminated)
		.almost_empty_data (),                                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                                      // (terminated)
		.out_empty         (),                                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                                      // (terminated)
		.out_error         (),                                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                                      // (terminated)
		.out_channel       ()                                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) leds_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (leds_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (leds_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (leds_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (leds_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                              //                .channel
		.rf_sink_ready           (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                                                 //                .channel
		.rf_sink_ready           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) switches_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (switches_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switches_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switches_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switches_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switches_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switches_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switches_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switches_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switches_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switches_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switches_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switches_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switches_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switches_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                                 //                .channel
		.rf_sink_ready           (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) keys_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (keys_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (keys_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (keys_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (keys_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (keys_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (keys_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (keys_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (keys_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (keys_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (keys_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (keys_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (keys_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (keys_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (keys_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (keys_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (keys_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                             //                .channel
		.rf_sink_ready           (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                                   //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                                                   //       clk_reset.reset
		.m0_address              (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src13_ready),                                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src13_valid),                                                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_001_src13_data),                                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src13_startofpacket),                                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src13_endofpacket),                                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src13_channel),                                                                                     //                .channel
		.rf_sink_ready           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                                   //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                                                   // clk_reset.reset
		.in_data           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                                                 // (terminated)
		.csr_readdata      (),                                                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                                 // (terminated)
		.almost_full_data  (),                                                                                                                     // (terminated)
		.almost_empty_data (),                                                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                                                 // (terminated)
		.out_empty         (),                                                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                                                 // (terminated)
		.out_error         (),                                                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                                                 // (terminated)
		.out_channel       ()                                                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src14_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src14_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src14_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src14_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src14_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src14_channel),                                                              //                .channel
		.rf_sink_ready           (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ledr_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src15_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src15_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src15_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src15_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src15_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src15_channel),                                             //                .channel
		.rf_sink_ready           (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src16_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src16_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src16_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src16_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src16_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src16_channel),                                                            //                .channel
		.rf_sink_ready           (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) hex0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (hex0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src17_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src17_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src17_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src17_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src17_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src17_channel),                                             //                .channel
		.rf_sink_ready           (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) hex1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (hex1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src18_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src18_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src18_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src18_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src18_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src18_channel),                                             //                .channel
		.rf_sink_ready           (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) hex2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (hex2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src19_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src19_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src19_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src19_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src19_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src19_channel),                                             //                .channel
		.rf_sink_ready           (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) hex3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (hex3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src20_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src20_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src20_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src20_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src20_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src20_channel),                                             //                .channel
		.rf_sink_ready           (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (91),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) hex4_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (hex4_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex4_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex4_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex4_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex4_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex4_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex4_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src21_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src21_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src21_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src21_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src21_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src21_channel),                                             //                .channel
		.rf_sink_ready           (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (59),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (64),
		.PKT_SRC_ID_L              (60),
		.PKT_DEST_ID_H             (69),
		.PKT_DEST_ID_L             (65),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (73),
		.PKT_PROTECTION_L          (71),
		.PKT_RESPONSE_STATUS_H     (79),
		.PKT_RESPONSE_STATUS_L     (78),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (80),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                        //       clk_reset.reset
		.m0_address              (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_003_source0_ready),                                                                       //              cp.ready
		.cp_valid                (burst_adapter_003_source0_valid),                                                                       //                .valid
		.cp_data                 (burst_adapter_003_source0_data),                                                                        //                .data
		.cp_startofpacket        (burst_adapter_003_source0_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (burst_adapter_003_source0_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (burst_adapter_003_source0_channel),                                                                     //                .channel
		.rf_sink_ready           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (81),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                        // clk_reset.reset
		.in_data           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                                  // (terminated)
		.csr_readdata      (),                                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                  // (terminated)
		.almost_full_data  (),                                                                                                      // (terminated)
		.almost_empty_data (),                                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                                  // (terminated)
		.out_empty         (),                                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                                  // (terminated)
		.out_error         (),                                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                                  // (terminated)
		.out_channel       ()                                                                                                       // (terminated)
	);

	nios_system_addr_router addr_router (
		.sink_ready         (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                          //       src.ready
		.src_valid          (addr_router_src_valid),                                                                          //          .valid
		.src_data           (addr_router_src_data),                                                                           //          .data
		.src_channel        (addr_router_src_channel),                                                                        //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                     //          .endofpacket
	);

	nios_system_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                               //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                               //          .valid
		.src_data           (addr_router_001_src_data),                                                                //          .data
		.src_channel        (addr_router_001_src_channel),                                                             //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                          //          .endofpacket
	);

	nios_system_addr_router_002 addr_router_002 (
		.sink_ready         (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pixel_buffer_dma_0_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                         // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                                              //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                                              //          .valid
		.src_data           (addr_router_002_src_data),                                                                               //          .data
		.src_channel        (addr_router_002_src_channel),                                                                            //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                                      //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                                         //          .endofpacket
	);

	nios_system_id_router id_router (
		.sink_ready         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                          //       src.ready
		.src_valid          (id_router_src_valid),                                                                          //          .valid
		.src_data           (id_router_src_data),                                                                           //          .data
		.src_channel        (id_router_src_channel),                                                                        //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                     //          .endofpacket
	);

	nios_system_id_router_001 id_router_001 (
		.sink_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                             //       src.ready
		.src_valid          (id_router_001_src_valid),                                             //          .valid
		.src_data           (id_router_001_src_data),                                              //          .data
		.src_channel        (id_router_001_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                        //          .endofpacket
	);

	nios_system_id_router_002 id_router_002 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                //          .valid
		.src_data           (id_router_002_src_data),                                                                 //          .data
		.src_channel        (id_router_002_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                           //          .endofpacket
	);

	nios_system_id_router_002 id_router_003 (
		.sink_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                             //       src.ready
		.src_valid          (id_router_003_src_valid),                                             //          .valid
		.src_data           (id_router_003_src_data),                                              //          .data
		.src_channel        (id_router_003_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                        //          .endofpacket
	);

	nios_system_id_router_002 id_router_004 (
		.sink_ready         (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                 //       src.ready
		.src_valid          (id_router_004_src_valid),                                                 //          .valid
		.src_data           (id_router_004_src_data),                                                  //          .data
		.src_channel        (id_router_004_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                            //          .endofpacket
	);

	nios_system_id_router_005 id_router_005 (
		.sink_ready         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                   //          .valid
		.src_data           (id_router_005_src_data),                                                                    //          .data
		.src_channel        (id_router_005_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                              //          .endofpacket
	);

	nios_system_id_router_002 id_router_006 (
		.sink_ready         (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pixel_buffer_dma_0_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                            //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                            //          .valid
		.src_data           (id_router_006_src_data),                                                                             //          .data
		.src_channel        (id_router_006_src_channel),                                                                          //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                                    //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                                       //          .endofpacket
	);

	nios_system_id_router_002 id_router_007 (
		.sink_ready         (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                                          //       src.ready
		.src_valid          (id_router_007_src_valid),                                                                          //          .valid
		.src_data           (id_router_007_src_data),                                                                           //          .data
		.src_channel        (id_router_007_src_channel),                                                                        //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                                     //          .endofpacket
	);

	nios_system_id_router_008 id_router_008 (
		.sink_ready         (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                         //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                         //          .valid
		.src_data           (id_router_008_src_data),                                                                          //          .data
		.src_channel        (id_router_008_src_channel),                                                                       //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                                 //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                                    //          .endofpacket
	);

	nios_system_id_router_002 id_router_009 (
		.sink_ready         (leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (leds_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                            //       src.ready
		.src_valid          (id_router_009_src_valid),                                            //          .valid
		.src_data           (id_router_009_src_data),                                             //          .data
		.src_channel        (id_router_009_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                       //          .endofpacket
	);

	nios_system_id_router_002 id_router_010 (
		.sink_ready         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                                //       src.ready
		.src_valid          (id_router_010_src_valid),                                                                //          .valid
		.src_data           (id_router_010_src_data),                                                                 //          .data
		.src_channel        (id_router_010_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                           //          .endofpacket
	);

	nios_system_id_router_002 id_router_011 (
		.sink_ready         (switches_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switches_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switches_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switches_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                //       src.ready
		.src_valid          (id_router_011_src_valid),                                                //          .valid
		.src_data           (id_router_011_src_data),                                                 //          .data
		.src_channel        (id_router_011_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                           //          .endofpacket
	);

	nios_system_id_router_002 id_router_012 (
		.sink_ready         (keys_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (keys_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (keys_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (keys_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (keys_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                            //       src.ready
		.src_valid          (id_router_012_src_valid),                                            //          .valid
		.src_data           (id_router_012_src_data),                                             //          .data
		.src_channel        (id_router_012_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                       //          .endofpacket
	);

	nios_system_id_router_002 id_router_013 (
		.sink_ready         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                                         //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                                         // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                                                    //       src.ready
		.src_valid          (id_router_013_src_valid),                                                                                    //          .valid
		.src_data           (id_router_013_src_data),                                                                                     //          .data
		.src_channel        (id_router_013_src_channel),                                                                                  //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                                                            //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                                                               //          .endofpacket
	);

	nios_system_id_router_002 id_router_014 (
		.sink_ready         (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                             //       src.ready
		.src_valid          (id_router_014_src_valid),                                                             //          .valid
		.src_data           (id_router_014_src_data),                                                              //          .data
		.src_channel        (id_router_014_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                                        //          .endofpacket
	);

	nios_system_id_router_002 id_router_015 (
		.sink_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                            //       src.ready
		.src_valid          (id_router_015_src_valid),                                            //          .valid
		.src_data           (id_router_015_src_data),                                             //          .data
		.src_channel        (id_router_015_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                       //          .endofpacket
	);

	nios_system_id_router_002 id_router_016 (
		.sink_ready         (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                           //       src.ready
		.src_valid          (id_router_016_src_valid),                                                           //          .valid
		.src_data           (id_router_016_src_data),                                                            //          .data
		.src_channel        (id_router_016_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                                      //          .endofpacket
	);

	nios_system_id_router_002 id_router_017 (
		.sink_ready         (hex0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                            //       src.ready
		.src_valid          (id_router_017_src_valid),                                            //          .valid
		.src_data           (id_router_017_src_data),                                             //          .data
		.src_channel        (id_router_017_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                       //          .endofpacket
	);

	nios_system_id_router_002 id_router_018 (
		.sink_ready         (hex1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                            //       src.ready
		.src_valid          (id_router_018_src_valid),                                            //          .valid
		.src_data           (id_router_018_src_data),                                             //          .data
		.src_channel        (id_router_018_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                       //          .endofpacket
	);

	nios_system_id_router_002 id_router_019 (
		.sink_ready         (hex2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                            //       src.ready
		.src_valid          (id_router_019_src_valid),                                            //          .valid
		.src_data           (id_router_019_src_data),                                             //          .data
		.src_channel        (id_router_019_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                       //          .endofpacket
	);

	nios_system_id_router_002 id_router_020 (
		.sink_ready         (hex3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                            //       src.ready
		.src_valid          (id_router_020_src_valid),                                            //          .valid
		.src_data           (id_router_020_src_data),                                             //          .data
		.src_channel        (id_router_020_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                       //          .endofpacket
	);

	nios_system_id_router_002 id_router_021 (
		.sink_ready         (hex4_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex4_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex4_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                            //       src.ready
		.src_valid          (id_router_021_src_valid),                                            //          .valid
		.src_data           (id_router_021_src_data),                                             //          .data
		.src_channel        (id_router_021_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                       //          .endofpacket
	);

	nios_system_id_router_008 id_router_022 (
		.sink_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_022_src_valid),                                                                     //          .valid
		.src_data           (id_router_022_src_data),                                                                      //          .data
		.src_channel        (id_router_022_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)                                                                //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (23),
		.VALID_WIDTH               (23),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clocks_sys_clk_clk),             //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (92),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (23),
		.VALID_WIDTH               (23),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clocks_sys_clk_clk),                 //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (68),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (23),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (clocks_sys_clk_clk),                  //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_001_src_valid),          //     sink0.valid
		.sink0_data            (cmd_xbar_mux_001_src_data),           //          .data
		.sink0_channel         (cmd_xbar_mux_001_src_channel),        //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_001_src_startofpacket),  //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_001_src_endofpacket),    //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_001_src_ready),          //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (68),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (23),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_001 (
		.clk                   (clocks_sys_clk_clk),                      //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_005_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_005_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_005_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_005_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_005_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_005_src_ready),              //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (59),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (80),
		.ST_CHANNEL_W              (23),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_002 (
		.clk                   (clocks_sys_clk_clk),                      //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_003_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_003_src_data),              //          .data
		.sink0_channel         (width_adapter_003_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_003_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_003_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_003_src_ready),             //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (59),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (80),
		.ST_CHANNEL_W              (23),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_003 (
		.clk                   (clocks_sys_clk_clk),                      //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_004_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_004_src_data),              //          .data
		.sink0_channel         (width_adapter_004_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_004_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_004_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_004_src_ready),             //          .ready
		.source0_valid         (burst_adapter_003_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_003_source0_data),          //          .data
		.source0_channel       (burst_adapter_003_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_003_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_003_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_003_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                                // reset_in0.reset
		.reset_in1  (nios2_processor_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clocks_sys_clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),                // reset_out.reset
		.reset_in2  (1'b0),                                          // (terminated)
		.reset_in3  (1'b0),                                          // (terminated)
		.reset_in4  (1'b0),                                          // (terminated)
		.reset_in5  (1'b0),                                          // (terminated)
		.reset_in6  (1'b0),                                          // (terminated)
		.reset_in7  (1'b0),                                          // (terminated)
		.reset_in8  (1'b0),                                          // (terminated)
		.reset_in9  (1'b0),                                          // (terminated)
		.reset_in10 (1'b0),                                          // (terminated)
		.reset_in11 (1'b0),                                          // (terminated)
		.reset_in12 (1'b0),                                          // (terminated)
		.reset_in13 (1'b0),                                          // (terminated)
		.reset_in14 (1'b0),                                          // (terminated)
		.reset_in15 (1'b0)                                           // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                                // reset_in0.reset
		.reset_in1  (nios2_processor_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                                       //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),            // reset_out.reset
		.reset_in2  (1'b0),                                          // (terminated)
		.reset_in3  (1'b0),                                          // (terminated)
		.reset_in4  (1'b0),                                          // (terminated)
		.reset_in5  (1'b0),                                          // (terminated)
		.reset_in6  (1'b0),                                          // (terminated)
		.reset_in7  (1'b0),                                          // (terminated)
		.reset_in8  (1'b0),                                          // (terminated)
		.reset_in9  (1'b0),                                          // (terminated)
		.reset_in10 (1'b0),                                          // (terminated)
		.reset_in11 (1'b0),                                          // (terminated)
		.reset_in12 (1'b0),                                          // (terminated)
		.reset_in13 (1'b0),                                          // (terminated)
		.reset_in14 (1'b0),                                          // (terminated)
		.reset_in15 (1'b0)                                           // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (nios2_processor_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                                // reset_in1.reset
		.clk        (clocks_vga_clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset),            // reset_out.reset
		.reset_in2  (1'b0),                                          // (terminated)
		.reset_in3  (1'b0),                                          // (terminated)
		.reset_in4  (1'b0),                                          // (terminated)
		.reset_in5  (1'b0),                                          // (terminated)
		.reset_in6  (1'b0),                                          // (terminated)
		.reset_in7  (1'b0),                                          // (terminated)
		.reset_in8  (1'b0),                                          // (terminated)
		.reset_in9  (1'b0),                                          // (terminated)
		.reset_in10 (1'b0),                                          // (terminated)
		.reset_in11 (1'b0),                                          // (terminated)
		.reset_in12 (1'b0),                                          // (terminated)
		.reset_in13 (1'b0),                                          // (terminated)
		.reset_in14 (1'b0),                                          // (terminated)
		.reset_in15 (1'b0)                                           // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_003 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clocks_sys_clk_clk),                 //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clocks_sys_clk_clk),                //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //           .endofpacket
	);

	nios_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clocks_sys_clk_clk),                     //        clk.clk
		.reset               (rst_controller_reset_out_reset),         //  clk_reset.reset
		.sink_ready          (limiter_001_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_001_cmd_src_channel),            //           .channel
		.sink_data           (limiter_001_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_001_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_001_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_001_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //           .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //      src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //           .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //           .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //           .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //           .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //           .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //      src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //           .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //           .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //           .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //           .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //           .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //      src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //           .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //           .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //           .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //           .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket),   //           .endofpacket
		.src17_ready         (cmd_xbar_demux_001_src17_ready),         //      src17.ready
		.src17_valid         (cmd_xbar_demux_001_src17_valid),         //           .valid
		.src17_data          (cmd_xbar_demux_001_src17_data),          //           .data
		.src17_channel       (cmd_xbar_demux_001_src17_channel),       //           .channel
		.src17_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //           .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_001_src17_endofpacket),   //           .endofpacket
		.src18_ready         (cmd_xbar_demux_001_src18_ready),         //      src18.ready
		.src18_valid         (cmd_xbar_demux_001_src18_valid),         //           .valid
		.src18_data          (cmd_xbar_demux_001_src18_data),          //           .data
		.src18_channel       (cmd_xbar_demux_001_src18_channel),       //           .channel
		.src18_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //           .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_001_src18_endofpacket),   //           .endofpacket
		.src19_ready         (cmd_xbar_demux_001_src19_ready),         //      src19.ready
		.src19_valid         (cmd_xbar_demux_001_src19_valid),         //           .valid
		.src19_data          (cmd_xbar_demux_001_src19_data),          //           .data
		.src19_channel       (cmd_xbar_demux_001_src19_channel),       //           .channel
		.src19_startofpacket (cmd_xbar_demux_001_src19_startofpacket), //           .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_001_src19_endofpacket),   //           .endofpacket
		.src20_ready         (cmd_xbar_demux_001_src20_ready),         //      src20.ready
		.src20_valid         (cmd_xbar_demux_001_src20_valid),         //           .valid
		.src20_data          (cmd_xbar_demux_001_src20_data),          //           .data
		.src20_channel       (cmd_xbar_demux_001_src20_channel),       //           .channel
		.src20_startofpacket (cmd_xbar_demux_001_src20_startofpacket), //           .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_001_src20_endofpacket),   //           .endofpacket
		.src21_ready         (cmd_xbar_demux_001_src21_ready),         //      src21.ready
		.src21_valid         (cmd_xbar_demux_001_src21_valid),         //           .valid
		.src21_data          (cmd_xbar_demux_001_src21_data),          //           .data
		.src21_channel       (cmd_xbar_demux_001_src21_channel),       //           .channel
		.src21_startofpacket (cmd_xbar_demux_001_src21_startofpacket), //           .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_001_src21_endofpacket),   //           .endofpacket
		.src22_ready         (cmd_xbar_demux_001_src22_ready),         //      src22.ready
		.src22_valid         (cmd_xbar_demux_001_src22_valid),         //           .valid
		.src22_data          (cmd_xbar_demux_001_src22_data),          //           .data
		.src22_channel       (cmd_xbar_demux_001_src22_channel),       //           .channel
		.src22_startofpacket (cmd_xbar_demux_001_src22_startofpacket), //           .startofpacket
		.src22_endofpacket   (cmd_xbar_demux_001_src22_endofpacket)    //           .endofpacket
	);

	nios_system_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux_001 cmd_xbar_mux_001 (
		.clk                 (clocks_sys_clk_clk),                  //       clk.clk
		.reset               (rst_controller_reset_out_reset),      // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),          //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),          //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),           //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),        //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),  //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),    //          .endofpacket
		.sink0_ready         (width_adapter_src_ready),             //     sink0.ready
		.sink0_valid         (width_adapter_src_valid),             //          .valid
		.sink0_channel       (width_adapter_src_channel),           //          .channel
		.sink0_data          (width_adapter_src_data),              //          .data
		.sink0_startofpacket (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (width_adapter_src_endofpacket),       //          .endofpacket
		.sink1_ready         (width_adapter_001_src_ready),         //     sink1.ready
		.sink1_valid         (width_adapter_001_src_valid),         //          .valid
		.sink1_channel       (width_adapter_001_src_channel),       //          .channel
		.sink1_data          (width_adapter_001_src_data),          //          .data
		.sink1_startofpacket (width_adapter_001_src_startofpacket), //          .startofpacket
		.sink1_endofpacket   (width_adapter_001_src_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux_001 cmd_xbar_mux_005 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_002_src_ready),           //     sink0.ready
		.sink0_valid         (width_adapter_002_src_valid),           //          .valid
		.sink0_channel       (width_adapter_002_src_channel),         //          .channel
		.sink0_data          (width_adapter_002_src_data),            //          .data
		.sink0_startofpacket (width_adapter_002_src_startofpacket),   //          .startofpacket
		.sink0_endofpacket   (width_adapter_002_src_endofpacket),     //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clocks_sys_clk_clk),                //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_005 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_006 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_007 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_008 rsp_xbar_demux_008 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_009 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_010 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_011 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_012 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_013 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_014 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_015 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_016 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_017 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_018 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_019 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_020 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_021 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_021_src_ready),               //      sink.ready
		.sink_channel       (id_router_021_src_channel),             //          .channel
		.sink_data          (id_router_021_src_data),                //          .data
		.sink_startofpacket (id_router_021_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_021_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_021_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_008 rsp_xbar_demux_022 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_022_src_ready),               //      sink.ready
		.sink_channel       (id_router_022_src_channel),             //          .channel
		.sink_data          (id_router_022_src_data),                //          .data
		.sink_startofpacket (id_router_022_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_022_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_022_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clocks_sys_clk_clk),                  //       clk.clk
		.reset               (rst_controller_reset_out_reset),      // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),              //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),              //          .valid
		.src_data            (rsp_xbar_mux_src_data),               //          .data
		.src_channel         (rsp_xbar_mux_src_channel),            //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),      //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),        //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),           //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),           //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),         //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),            //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),   //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),     //          .endofpacket
		.sink1_ready         (width_adapter_005_src_ready),         //     sink1.ready
		.sink1_valid         (width_adapter_005_src_valid),         //          .valid
		.sink1_channel       (width_adapter_005_src_channel),       //          .channel
		.sink1_data          (width_adapter_005_src_data),          //          .data
		.sink1_startofpacket (width_adapter_005_src_startofpacket), //          .startofpacket
		.sink1_endofpacket   (width_adapter_005_src_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (width_adapter_006_src_ready),           //     sink1.ready
		.sink1_valid          (width_adapter_006_src_valid),           //          .valid
		.sink1_channel        (width_adapter_006_src_channel),         //          .channel
		.sink1_data           (width_adapter_006_src_data),            //          .data
		.sink1_startofpacket  (width_adapter_006_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket    (width_adapter_006_src_endofpacket),     //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (width_adapter_007_src_ready),           //     sink5.ready
		.sink5_valid          (width_adapter_007_src_valid),           //          .valid
		.sink5_channel        (width_adapter_007_src_channel),         //          .channel
		.sink5_data           (width_adapter_007_src_data),            //          .data
		.sink5_startofpacket  (width_adapter_007_src_startofpacket),   //          .startofpacket
		.sink5_endofpacket    (width_adapter_007_src_endofpacket),     //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (width_adapter_008_src_ready),           //     sink8.ready
		.sink8_valid          (width_adapter_008_src_valid),           //          .valid
		.sink8_channel        (width_adapter_008_src_channel),         //          .channel
		.sink8_data           (width_adapter_008_src_data),            //          .data
		.sink8_startofpacket  (width_adapter_008_src_startofpacket),   //          .startofpacket
		.sink8_endofpacket    (width_adapter_008_src_endofpacket),     //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_019_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_020_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.sink21_ready         (rsp_xbar_demux_021_src0_ready),         //    sink21.ready
		.sink21_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.sink21_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.sink21_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.sink21_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.sink21_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.sink22_ready         (width_adapter_009_src_ready),           //    sink22.ready
		.sink22_valid         (width_adapter_009_src_valid),           //          .valid
		.sink22_channel       (width_adapter_009_src_channel),         //          .channel
		.sink22_data          (width_adapter_009_src_data),            //          .data
		.sink22_startofpacket (width_adapter_009_src_startofpacket),   //          .startofpacket
		.sink22_endofpacket   (width_adapter_009_src_endofpacket)      //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (88),
		.OUT_PKT_RESPONSE_STATUS_L     (87),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (23),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (clocks_sys_clk_clk),                //       clk.clk
		.reset                (rst_controller_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src1_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_src1_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_src1_ready),         //          .ready
		.in_data              (cmd_xbar_demux_src1_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_src_data),            //          .data
		.out_channel          (width_adapter_src_channel),         //          .channel
		.out_valid            (width_adapter_src_valid),           //          .valid
		.out_ready            (width_adapter_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                             // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (88),
		.OUT_PKT_RESPONSE_STATUS_L     (87),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (23),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_001 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src1_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src1_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src1_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src1_data),          //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_001_src_data),            //          .data
		.out_channel          (width_adapter_001_src_channel),         //          .channel
		.out_valid            (width_adapter_001_src_valid),           //          .valid
		.out_ready            (width_adapter_001_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (88),
		.OUT_PKT_RESPONSE_STATUS_L     (87),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (23),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_002 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src5_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src5_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src5_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src5_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src5_data),          //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_002_src_data),            //          .data
		.out_channel          (width_adapter_002_src_channel),         //          .channel
		.out_valid            (width_adapter_002_src_valid),           //          .valid
		.out_ready            (width_adapter_002_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (79),
		.OUT_PKT_RESPONSE_STATUS_L     (78),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (80),
		.ST_CHANNEL_W                  (23),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_003 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src8_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src8_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src8_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src8_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src8_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src8_data),          //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_003_src_data),            //          .data
		.out_channel          (width_adapter_003_src_channel),         //          .channel
		.out_valid            (width_adapter_003_src_valid),           //          .valid
		.out_ready            (width_adapter_003_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (79),
		.OUT_PKT_RESPONSE_STATUS_L     (78),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (80),
		.ST_CHANNEL_W                  (23),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_004 (
		.clk                  (clocks_sys_clk_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src22_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src22_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src22_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src22_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src22_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src22_data),          //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_004_src_data),             //          .data
		.out_channel          (width_adapter_004_src_channel),          //          .channel
		.out_valid            (width_adapter_004_src_valid),            //          .valid
		.out_ready            (width_adapter_004_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (88),
		.IN_PKT_RESPONSE_STATUS_L      (87),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (23),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_005 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_001_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_001_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_001_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_001_src0_data),          //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_005_src_data),            //          .data
		.out_channel          (width_adapter_005_src_channel),         //          .channel
		.out_valid            (width_adapter_005_src_valid),           //          .valid
		.out_ready            (width_adapter_005_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (88),
		.IN_PKT_RESPONSE_STATUS_L      (87),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (23),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_006 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_001_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_001_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_001_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_001_src1_data),          //          .data
		.out_endofpacket      (width_adapter_006_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_006_src_data),            //          .data
		.out_channel          (width_adapter_006_src_channel),         //          .channel
		.out_valid            (width_adapter_006_src_valid),           //          .valid
		.out_ready            (width_adapter_006_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_006_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (88),
		.IN_PKT_RESPONSE_STATUS_L      (87),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (23),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_007 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_005_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_005_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_005_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_005_src0_data),          //          .data
		.out_endofpacket      (width_adapter_007_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_007_src_data),            //          .data
		.out_channel          (width_adapter_007_src_channel),         //          .channel
		.out_valid            (width_adapter_007_src_valid),           //          .valid
		.out_ready            (width_adapter_007_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_007_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (79),
		.IN_PKT_RESPONSE_STATUS_L      (78),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (80),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (23),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_008 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_008_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_008_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_008_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_008_src0_data),          //          .data
		.out_endofpacket      (width_adapter_008_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_008_src_data),            //          .data
		.out_channel          (width_adapter_008_src_channel),         //          .channel
		.out_valid            (width_adapter_008_src_valid),           //          .valid
		.out_ready            (width_adapter_008_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_008_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (79),
		.IN_PKT_RESPONSE_STATUS_L      (78),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (80),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (23),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_009 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_022_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_022_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_022_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_022_src0_data),          //          .data
		.out_endofpacket      (width_adapter_009_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_009_src_data),            //          .data
		.out_channel          (width_adapter_009_src_channel),         //          .channel
		.out_valid            (width_adapter_009_src_valid),           //          .valid
		.out_ready            (width_adapter_009_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_009_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clocks_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.sender_irq    (nios2_processor_d_irq_irq)       //    sender.irq
	);

endmodule
